///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_RV32ZBA
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_rv32zba_t;


covergroup sh1add_cg with function sample(ins_rv32zba_t ins);
    option.per_instance = 1; 
    option.comment = "sh1add";
    cp_asm_count : coverpoint ins.ins_str == "sh1add"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  =    {0};
        wildcard bins one  =     {32'b00000000000000000000000000000001};
        wildcard bins two  =     {32'b00000000000000000000000000000010};
        wildcard bins min  =     {32'b10000000000000000000000000000000};
        wildcard bins minp1  =   {32'b10000000000000000000000000000001};
        wildcard bins max  =     {32'b01111111111111111111111111111111};
        wildcard bins maxm1  =   {32'b01111111111111111111111111111110};
        wildcard bins ones  =    {32'b11111111111111111111111111111111};
        wildcard bins onesm1  =  {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
endgroup

covergroup sh2add_cg with function sample(ins_rv32zba_t ins);
    option.per_instance = 1; 
    option.comment = "sh2add";
    cp_asm_count : coverpoint ins.ins_str == "sh2add"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  =    {0};
        wildcard bins one  =     {32'b00000000000000000000000000000001};
        wildcard bins two  =     {32'b00000000000000000000000000000010};
        wildcard bins min  =     {32'b10000000000000000000000000000000};
        wildcard bins minp1  =   {32'b10000000000000000000000000000001};
        wildcard bins max  =     {32'b01111111111111111111111111111111};
        wildcard bins maxm1  =   {32'b01111111111111111111111111111110};
        wildcard bins ones  =    {32'b11111111111111111111111111111111};
        wildcard bins onesm1  =  {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
endgroup

covergroup sh3add_cg with function sample(ins_rv32zba_t ins);
    option.per_instance = 1; 
    option.comment = "sh3add";
    cp_asm_count : coverpoint ins.ins_str == "sh3add"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  =    {0};
        wildcard bins one  =     {32'b00000000000000000000000000000001};
        wildcard bins two  =     {32'b00000000000000000000000000000010};
        wildcard bins min  =     {32'b10000000000000000000000000000000};
        wildcard bins minp1  =   {32'b10000000000000000000000000000001};
        wildcard bins max  =     {32'b01111111111111111111111111111111};
        wildcard bins maxm1  =   {32'b01111111111111111111111111111110};
        wildcard bins ones  =    {32'b11111111111111111111111111111111};
        wildcard bins onesm1  =  {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one  = {32'b00000000000000000000000000000001};
        wildcard bins two  = {32'b00000000000000000000000000000010};
        wildcard bins min  = {32'b10000000000000000000000000000000};
        wildcard bins minp1  = {32'b10000000000000000000000000000001};
        wildcard bins max  = {32'b01111111111111111111111111111111};
        wildcard bins maxm1  = {32'b01111111111111111111111111111110};
        wildcard bins ones  = {32'b11111111111111111111111111111111};
        wildcard bins onesm1  = {32'b11111111111111111111111111111110};
        wildcard bins walkeodd = {32'b10101010101010101010101010101010};
        wildcard bins walkeven = {32'b01010101010101010101010101010101};
        wildcard bins random   = {32'b01011011101111001000100001110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
endgroup

function void rv32zba_sample(int hart, int issue);
    ins_rv32zba_t ins;

    case (traceDataQ[hart][issue][0].inst_name)
        "sh1add"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sh1add_cg.sample(ins); 
        end
        "sh2add"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sh2add_cg.sample(ins); 
        end
        "sh3add"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sh3add_cg.sample(ins); 
        end
    endcase
endfunction
