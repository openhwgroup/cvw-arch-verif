///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    amoadd_w_cg = new(); amoadd_w_cg.set_inst_name("obj_amoadd_w");
    amoand_w_cg = new(); amoand_w_cg.set_inst_name("obj_amoand_w");
    amoaxor_w_cg = new(); amoaxor_w_cg.set_inst_name("obj_amoaxor_w");
    amomax_w_cg = new(); amomax_w_cg.set_inst_name("obj_amomax_w");
    amomaxu_w_cg = new(); amomaxu_w_cg.set_inst_name("obj_amomaxu_w");
    amomin_w_cg = new(); amomin_w_cg.set_inst_name("obj_amomin_w");
    amominu_w_cg = new(); amominu_w_cg.set_inst_name("obj_amominu_w");
    amoor_w_cg = new(); amoor_w_cg.set_inst_name("obj_amoor_w");
    amoswap_w_cg = new(); amoswap_w_cg.set_inst_name("obj_amoswap_w");
