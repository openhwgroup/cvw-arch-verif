///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fadd_d_cg = new(); fadd_d_cg.set_inst_name("obj_fadd_d");
    fclass_d_cg = new(); fclass_d_cg.set_inst_name("obj_fclass_d");
    fcvt_d_l_cg = new(); fcvt_d_l_cg.set_inst_name("obj_fcvt_d_l");
    fcvt_d_lu_cg = new(); fcvt_d_lu_cg.set_inst_name("obj_fcvt_d_lu");
    fcvt_d_s_cg = new(); fcvt_d_s_cg.set_inst_name("obj_fcvt_d_s");
    fcvt_d_w_cg = new(); fcvt_d_w_cg.set_inst_name("obj_fcvt_d_w");
    fcvt_d_wu_cg = new(); fcvt_d_wu_cg.set_inst_name("obj_fcvt_d_wu");
    fcvt_l_d_cg = new(); fcvt_l_d_cg.set_inst_name("obj_fcvt_l_d");
    fcvt_lu_d_cg = new(); fcvt_lu_d_cg.set_inst_name("obj_fcvt_lu_d");
    fcvt_s_d_cg = new(); fcvt_s_d_cg.set_inst_name("obj_fcvt_s_d");
    fcvt_w_d_cg = new(); fcvt_w_d_cg.set_inst_name("obj_fcvt_w_d");
    fcvt_wu_d_cg = new(); fcvt_wu_d_cg.set_inst_name("obj_fcvt_wu_d");
    fdiv_d_cg = new(); fdiv_d_cg.set_inst_name("obj_fdiv_d");
    feq_d_cg = new(); feq_d_cg.set_inst_name("obj_feq_d");
    fld_cg = new(); fld_cg.set_inst_name("obj_fld");
    fle_d_cg = new(); fle_d_cg.set_inst_name("obj_fle_d");
    flt_d_cg = new(); flt_d_cg.set_inst_name("obj_flt_d");
    fmadd_d_cg = new(); fmadd_d_cg.set_inst_name("obj_fmadd_d");
    fmax_d_cg = new(); fmax_d_cg.set_inst_name("obj_fmax_d");
    fmin_d_cg = new(); fmin_d_cg.set_inst_name("obj_fmin_d");
    fmsub_d_cg = new(); fmsub_d_cg.set_inst_name("obj_fmsub_d");
    fmul_d_cg = new(); fmul_d_cg.set_inst_name("obj_fmul_d");
    fmv_d_x_cg = new(); fmv_d_x_cg.set_inst_name("obj_fmv_d_x");
    fmv_x_d_cg = new(); fmv_x_d_cg.set_inst_name("obj_fmv_x_d");
    fnmadd_d_cg = new(); fnmadd_d_cg.set_inst_name("obj_fnmadd_d");
    fnmsub_d_cg = new(); fnmsub_d_cg.set_inst_name("obj_fnmsub_d");
    fsd_cg = new(); fsd_cg.set_inst_name("obj_fsd");
    fsgnj_d_cg = new(); fsgnj_d_cg.set_inst_name("obj_fsgnj_d");
    fsgnjn_d_cg = new(); fsgnjn_d_cg.set_inst_name("obj_fsgnjn_d");
    fsgnjx_d_cg = new(); fsgnjx_d_cg.set_inst_name("obj_fsgnjx_d");
    fsqrt_d_cg = new(); fsqrt_d_cg.set_inst_name("obj_fsqrt_d");
    fsub_d_cg = new(); fsub_d_cg.set_inst_name("obj_fsub_d");
