///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    lr_w_cg = new(); lr_w_cg.set_inst_name("obj_lr_w");
    sc_w_cg = new(); sc_w_cg.set_inst_name("obj_sc_w");
