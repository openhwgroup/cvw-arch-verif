///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ucsr_cg = new();         ucsr_cg.set_inst_name("obj_ucsr");
    uprivinst_cg = new();    uprivinst_cg.set_inst_name("obj_uprivinst");
