///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    SsstrictM_instr_cg = new();        SsstrictM_instr_cg.set_inst_name("obj_SsstrictM_instr");
    SsstrictM_comp_instr_cg = new();   SsstrictM_comp_instr_cg.set_inst_name("obj_SsstrictM_comp_instr");
     
