    `include "RV64VM_coverage.svh"
    `include "RV64VM_PMP_coverage.svh"
    `include "RV64Zicbom_coverage.svh"
