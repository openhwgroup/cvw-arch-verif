///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    RV64VM_satp_cg = new(); RV64VM_satp_cg.set_inst_name("obj_RV64VM_satp");
    RV64VM_PA_VA_cg = new(); RV64VM_PA_VA_cg.set_inst_name("obj_RV64VM_PA_VA");
    RV64VM_sfence_cg = new(); RV64VM_sfence_cg.set_inst_name("obj_RV64VM_sfence");
    RV64VM_mstatus_mprv_cg = new(); RV64VM_mstatus_mprv_cg.set_inst_name("obj_RV64VM_mstatus_mprv");
    RV64VM_vm_permissions_cg = new(); RV64VM_vm_permissions_cg.set_inst_name("obj_RV64VM_vm_permissions");
    RV64VM_res_global_pte_cg = new(); RV64VM_res_global_pte_cg.set_inst_name("obj_RV64VM_res_global_pte");
    RV64VM_add_feature_cg = new(); RV64VM_add_feature_cg.set_inst_name("obj_RV64VM_add_feature");
