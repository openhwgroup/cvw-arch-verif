///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Standard Covergroups
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define RAMBASEADDR 32'h80000000
`define LARGESTPROGRAM 32'h00010000
`define SAFEREGIONSTART (`RAMBASEADDR + `LARGESTPROGRAM)
`define REGIONSTART `SAFEREGIONSTART
`define G 0
`define g (2**(max(`G,1)+2))
`define STANDARD_REGION (`REGIONSTART >> (`G+2)) | ((1 << (`G-1)) - 1)

`define COVER_RV32PMP
`define COVER_RV64PMP

covergroup PMPM_cg with function sample(ins_t ins, logic [XLEN-1:0] pmpcfg [3:0],  logic [XLEN-1:0] pmpaddr [14:0], logic [29:0] pmpcfg_rw, logic [29:0] pmpcfg_a, logic [14:0] pmpcfg_x, logic [14:0] pmpcfg_l, logic [14:0] pmp_hit);
    option.per_instance = 0;
    `include  "coverage/RISCV_coverage_standard_coverpoints.svh"

    addr_in_region: coverpoint (ins.current.rs1_val + ins.current.imm) {
        bins at_region     = {`REGIONSTART};
    }

    standard_region: coverpoint pmpaddr[0] {
        bins standard_region = {`STANDARD_REGION};
    }

    Mcause: coverpoint ins.current.csr[12'h342]{  
        bins illegal_ins  = {32'd2};
        bins no_exception = {32'd0};
    }

	locked_region: coverpoint pmpcfg_l[1] {
		bins locked = {1'b1};
	}
	
	unlocked_region: coverpoint pmpcfg_l[1] {
		bins unlocked = {1'b0};
	}
	
	pmpaddr_write_ignore: coverpoint (ins.current.csr[12'h3B1] == ins.prev.csr[12'h3B1]) {
		bins write_ignored  = {1};
	}

	pmpaddr_write_detect: coverpoint (ins.current.csr[12'h3B1] != ins.prev.csr[12'h3B1]) {
		bins write_detected  = {1};
	}

	pmpcfg_write_ignore: coverpoint (ins.current.csr[12'h3A1] == ins.prev.csr[12'h3A1]) {
		bins write_ignored  = {1};
	}

	pmpcfg_write_detect: coverpoint (ins.current.csr[12'h3A1] != ins.prev.csr[12'h3A1]) {
		bins write_detected  = {1};
	}

    pmp_region: coverpoint ins.current.csr[12'h3A0][12:11] {
        bins OFF   = {2'b00};
        bins TOR   = {2'b01};
        bins NAPOT = {2'b11};
    }

    exec_instr: coverpoint ins.current.insn {
        wildcard bins jalr = {32'b????????????_?????_000_?????_1100111};
    }

    read_instr: coverpoint ins.current.insn {
        wildcard bins lb  = {32'b????????????_?????_000_?????_0000011};
        wildcard bins lbu = {32'b????????????_?????_100_?????_0000011};
        wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
        wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
        wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
        `ifdef XLEN64
            wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
            wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
        `endif
    }

    write_instr: coverpoint ins.current.insn {
        wildcard bins sb = {32'b???????_?????_?????_000_?????_0100011};
        wildcard bins sh = {32'b???????_?????_?????_001_?????_0100011};
        wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
        `ifdef XLEN64
            wildcard bins sd = {32'b???????_?????_?????_011_?????_0100011};
        `endif
    }

    legal_lxwr: coverpoint pmpcfg[0][7:0] { 
            wildcard bins cfg_l000 = {8'b10011000};
            wildcard bins cfg_l001 = {8'b10011001};
            wildcard bins cfg_l011 = {8'b10011011};
            wildcard bins cfg_l100 = {8'b10011100};
            wildcard bins cfg_l101 = {8'b10011101};
            wildcard bins cfg_l111 = {8'b10011111};
    }
	
	X0: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 0, pmpcfg.L = 1 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_x0   = {75'b??????????????0_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_x0   = {75'b?????????????0?_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_x0   = {75'b????????????0??_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_x0   = {75'b???????????0???_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_x0   = {75'b??????????0????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_x0   = {75'b?????????0?????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_x0   = {75'b????????0??????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_x0   = {75'b???????0???????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_x0   = {75'b??????0????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_x0   = {75'b?????0?????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_x0  = {75'b????0??????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_x0  = {75'b???0???????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_x0  = {75'b??0????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_x0  = {75'b?0?????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_x0  = {75'b0??????????????_1??????????????_11????????????????????????????_1??????????????};
	}
	
	X1: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 1, pmpcfg.L = 1 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_x1   = {75'b??????????????1_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_x1   = {75'b?????????????1?_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_x1   = {75'b????????????1??_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_x1   = {75'b???????????1???_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_x1   = {75'b??????????1????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_x1   = {75'b?????????1?????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_x1   = {75'b????????1??????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_x1   = {75'b???????1???????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_x1   = {75'b??????1????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_x1   = {75'b?????1?????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_x1  = {75'b????1??????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_x1  = {75'b???1???????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_x1  = {75'b??1????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_x1  = {75'b?1?????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_x1  = {75'b1??????????????_1??????????????_11????????????????????????????_1??????????????};
	}
	
	RW00: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 0, pmpcfg.L = 1 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_rw00   = {90'b????????????????????????????00_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw00   = {90'b??????????????????????????00??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw00   = {90'b????????????????????????00????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw00   = {90'b??????????????????????00??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw00   = {90'b????????????????????00????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw00   = {90'b??????????????????00??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw00   = {90'b????????????????00????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw00   = {90'b??????????????00??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw00   = {90'b????????????00????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw00   = {90'b??????????00??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw00  = {90'b????????00????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw00  = {90'b??????00??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw00  = {90'b????00????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw00  = {90'b??00??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw00  = {90'b00????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}
	
	RW11: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 3, pmpcfg.L = 1 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????11_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????11??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????11????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????11??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????11????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????11??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????11????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????11??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw11     = {90'b????????????11????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw11     = {90'b??????????11??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw11    = {90'b????????11????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw11    = {90'b??????11??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw11    = {90'b????11????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw11    = {90'b??11??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw11    = {90'b11????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}
	
	RW10: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 1, pmpcfg.L = 1 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????01_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????01??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????01????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????01??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????01????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????01??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????01????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????01??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw11     = {90'b????????????01????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw11     = {90'b??????????01??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw11    = {90'b????????01????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw11    = {90'b??????01??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw11    = {90'b????01????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw11    = {90'b??01??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw11    = {90'b01????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}

	RWX000: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 0 and pmpcfg.A = 3 
		wildcard bins pmp0cfg_rwx000     = {105'b????????????????????????????00_??????????????0_??????????????0_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rwx000     = {105'b??????????????????????????00??_?????????????0?_?????????????0?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rwx000     = {105'b????????????????????????00????_????????????0??_????????????0??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rwx000     = {105'b??????????????????????00??????_???????????0???_???????????0???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rwx000     = {105'b????????????????????00????????_??????????0????_??????????0????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rwx000     = {105'b??????????????????00??????????_?????????0?????_?????????0?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rwx000     = {105'b????????????????00????????????_????????0??????_????????0??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rwx000     = {105'b??????????????00??????????????_???????0???????_???????0???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rwx000     = {105'b????????????00????????????????_??????0????????_??????0????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rwx000     = {105'b??????????00??????????????????_?????0?????????_?????0?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rwx000    = {105'b????????00????????????????????_????0??????????_????0??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rwx000    = {105'b??????00??????????????????????_???0???????????_???0???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rwx000    = {105'b????00????????????????????????_??0????????????_??0????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rwx000    = {105'b??00??????????????????????????_?0?????????????_?0?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rwx000    = {105'b00????????????????????????????_0??????????????_0??????????????_11????????????????????????????_1??????????????};
	}
	
    cp_cfg_X: cross priv_mode_m, legal_lxwr, exec_instr, standard_region, addr_in_region ;
    
    cp_cfg_R: cross priv_mode_m, legal_lxwr, read_instr, standard_region, addr_in_region ;

    cp_cfg_W: cross priv_mode_m, legal_lxwr, write_instr, standard_region, addr_in_region ;
	
	cp_cfg_X0_all: cross priv_mode_m, exec_instr, X0, addr_in_region ;
	
	cp_cfg_X1_all: cross priv_mode_m, exec_instr, X1, addr_in_region ;

	cp_cfg_Rw00_all: cross priv_mode_m, read_instr, RW00, addr_in_region ;

	cp_cfg_Rw10_all: cross priv_mode_m, read_instr, RW10, addr_in_region ;

	cp_cfg_Rw11_all: cross priv_mode_m, read_instr, RW11, addr_in_region ;

	cp_cfg_rW00_all: cross priv_mode_m, write_instr, RW00, addr_in_region ;

	cp_cfg_rW10_all: cross priv_mode_m, write_instr, RW10, addr_in_region ;

	cp_cfg_rW11_all: cross priv_mode_m, write_instr, RW11, addr_in_region ;

	cp_cfg_L_access_exec: cross priv_mode_m, exec_instr, RWX000, addr_in_region;

	cp_cfg_L_access_read: cross priv_mode_m, read_instr, RWX000, addr_in_region;

	cp_cfg_L_access_write: cross priv_mode_m, write_instr, RWX000, addr_in_region;

	cp_cfg_L1_pmpaddr: cross locked_region, pmp_region, pmpaddr_write_ignore; 

	cp_cfg_L0_pmpaddr: cross unlocked_region, pmp_region, pmpaddr_write_detect;

	cp_cfg_L1_pmpcfg: cross locked_region, pmp_region, pmpcfg_write_ignore; 

	cp_cfg_L0_pmpcfg: cross unlocked_region, pmp_region, pmpcfg_write_detect;
	
 
endgroup

function void pmp_sample(int hart, int issue, ins_t ins);

    logic [XLEN-1:0] pmpcfg [3:0];  
    logic [XLEN-1:0] pmpaddr [14:0]; 
    logic [29:0] pmpcfg_rw, pmpcfg_a;
    logic [14:0] pmpcfg_x, pmpcfg_l, pmp_hit;

    for (int i = 0; i < 4; i++) begin
        pmpcfg[i] = ins.current.csr[12'h3A0 + i];
    end
 
    for (int j = 0; j < 15; j++) begin
        pmpaddr[j] = ins.current.csr[12'h3B0 + j];
    end

	for (int k = 0; k < 15; k++) begin
	    pmp_hit[k] = (pmpaddr[k] == `STANDARD_REGION);
	end
	
	`ifdef XLEN32
		pmpcfg_rw = {
					 ins.current.csr[12'h3A3][17:16],
					 ins.current.csr[12'h3A3][9:8],
					 ins.current.csr[12'h3A3][1:0],
					 ins.current.csr[12'h3A2][25:24],
					 ins.current.csr[12'h3A2][17:16],
					 ins.current.csr[12'h3A2][9:8],
					 ins.current.csr[12'h3A2][1:0],
					 ins.current.csr[12'h3A1][25:24],
					 ins.current.csr[12'h3A1][17:16],
					 ins.current.csr[12'h3A1][9:8],
					 ins.current.csr[12'h3A1][1:0],
					 ins.current.csr[12'h3A0][25:24],
					 ins.current.csr[12'h3A0][17:16],
					 ins.current.csr[12'h3A0][9:8],
					 ins.current.csr[12'h3A0][1:0]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_rw = {
					 ins.current.csr[12'h3A2][49:48],
					 ins.current.csr[12'h3A2][41:40],
					 ins.current.csr[12'h3A2][33:32],
					 ins.current.csr[12'h3A2][25:24],
					 ins.current.csr[12'h3A2][17:16],
					 ins.current.csr[12'h3A2][9:8],
					 ins.current.csr[12'h3A2][1:0],
					 ins.current.csr[12'h3A0][57:56],
					 ins.current.csr[12'h3A0][49:48],
					 ins.current.csr[12'h3A0][41:40],
					 ins.current.csr[12'h3A0][33:32],
					 ins.current.csr[12'h3A0][25:24],
					 ins.current.csr[12'h3A0][17:16],
					 ins.current.csr[12'h3A0][9:8],
					 ins.current.csr[12'h3A0][1:0]
					};
	`endif
	
	`ifdef XLEN32
		pmpcfg_x =  {
					 ins.current.csr[12'h3A3][18],
					 ins.current.csr[12'h3A3][10],
					 ins.current.csr[12'h3A3][2],
					 ins.current.csr[12'h3A2][26],
					 ins.current.csr[12'h3A2][18],
					 ins.current.csr[12'h3A2][10],
					 ins.current.csr[12'h3A2][2],
					 ins.current.csr[12'h3A1][26],
					 ins.current.csr[12'h3A1][18],
					 ins.current.csr[12'h3A1][10],
					 ins.current.csr[12'h3A1][2],
					 ins.current.csr[12'h3A0][26],
					 ins.current.csr[12'h3A0][18],
					 ins.current.csr[12'h3A0][10],
					 ins.current.csr[12'h3A0][2]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_x =  {
					 ins.current.csr[12'h3A2][50],
					 ins.current.csr[12'h3A2][42],
					 ins.current.csr[12'h3A2][34],
					 ins.current.csr[12'h3A2][26],
					 ins.current.csr[12'h3A2][18],
					 ins.current.csr[12'h3A2][10],
					 ins.current.csr[12'h3A2][2],
					 ins.current.csr[12'h3A0][58],
					 ins.current.csr[12'h3A0][50],
					 ins.current.csr[12'h3A0][42],
					 ins.current.csr[12'h3A0][34],
					 ins.current.csr[12'h3A0][26],
					 ins.current.csr[12'h3A0][18],
					 ins.current.csr[12'h3A0][10],
					 ins.current.csr[12'h3A0][2]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_a =  {
					 ins.current.csr[12'h3A3][20:19],
					 ins.current.csr[12'h3A3][12:11],
					 ins.current.csr[12'h3A3][4:3],
					 ins.current.csr[12'h3A2][28:27],
					 ins.current.csr[12'h3A2][20:19],
					 ins.current.csr[12'h3A2][12:11],
					 ins.current.csr[12'h3A2][4:3],
					 ins.current.csr[12'h3A1][28:27],
					 ins.current.csr[12'h3A1][20:19],
					 ins.current.csr[12'h3A1][12:11],
					 ins.current.csr[12'h3A1][4:3],
					 ins.current.csr[12'h3A0][28:27],
					 ins.current.csr[12'h3A0][20:19],
					 ins.current.csr[12'h3A0][12:11],
					 ins.current.csr[12'h3A0][4:3]
					};
	`endif
	
	`ifdef XLEN64
		pmpcfg_a =  {
					 ins.current.csr[12'h3A2][52:51],
					 ins.current.csr[12'h3A2][44:43],
					 ins.current.csr[12'h3A2][36:35],
					 ins.current.csr[12'h3A2][28:27],
					 ins.current.csr[12'h3A2][20:19],
					 ins.current.csr[12'h3A2][12:11],
					 ins.current.csr[12'h3A2][4:3],
					 ins.current.csr[12'h3A0][60:59],
					 ins.current.csr[12'h3A0][52:51],
					 ins.current.csr[12'h3A0][44:43],
					 ins.current.csr[12'h3A0][36:35],
					 ins.current.csr[12'h3A0][28:27],
					 ins.current.csr[12'h3A0][20:19],
					 ins.current.csr[12'h3A0][12:11],
					 ins.current.csr[12'h3A0][4:3]
					};
	`endif
	
	`ifdef XLEN32
		pmpcfg_l =  {
					 ins.current.csr[12'h3A3][23],
					 ins.current.csr[12'h3A3][15],
					 ins.current.csr[12'h3A3][7],
					 ins.current.csr[12'h3A2][31],
					 ins.current.csr[12'h3A2][23],
					 ins.current.csr[12'h3A2][15],
					 ins.current.csr[12'h3A2][7],
					 ins.current.csr[12'h3A1][31],
					 ins.current.csr[12'h3A1][23],
					 ins.current.csr[12'h3A1][15],
					 ins.current.csr[12'h3A1][7],
					 ins.current.csr[12'h3A0][31],
					 ins.current.csr[12'h3A0][23],
					 ins.current.csr[12'h3A0][15],
					 ins.current.csr[12'h3A0][7]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_l =  {
					 ins.current.csr[12'h3A2][55],
					 ins.current.csr[12'h3A2][47],
					 ins.current.csr[12'h3A2][39],
					 ins.current.csr[12'h3A2][31],
					 ins.current.csr[12'h3A2][23],
					 ins.current.csr[12'h3A2][15],
					 ins.current.csr[12'h3A2][7],
					 ins.current.csr[12'h3A0][63],
					 ins.current.csr[12'h3A0][55],
					 ins.current.csr[12'h3A0][47],
					 ins.current.csr[12'h3A0][39],
					 ins.current.csr[12'h3A0][31],
					 ins.current.csr[12'h3A0][23],
					 ins.current.csr[12'h3A0][15],
					 ins.current.csr[12'h3A0][7]
					};
	`endif

    PMPM_cg.sample(ins, pmpcfg, pmpaddr, pmpcfg_rw, pmpcfg_a, pmpcfg_x, pmpcfg_l, pmp_hit); 
endfunction

