///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2025 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    SsstrictV_instr_cg = new();        SsstrictV_instr_cg.set_inst_name("obj_SsstrictV_instr");
    SsstrictV_vcsr_cg = new();         SsstrictV_vcsr_cg.set_inst_name("obj_SsstrictV_vcsr");
