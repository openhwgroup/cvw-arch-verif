///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    aes64esi_cg = new(); aes64esi_cg.set_inst_name("obj_aes64esi");
    aes64esmi_cg = new(); aes64esmi_cg.set_inst_name("obj_aes64esmi");
    aes64im_cg = new(); aes64im_cg.set_inst_name("obj_aes64im");
    aes64ks1i_cg = new(); aes64ks1i_cg.set_inst_name("obj_aes64ks1i");
    aes64ks2_cg = new(); aes64ks2_cg.set_inst_name("obj_aes64ks2");
