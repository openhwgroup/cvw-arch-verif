///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Standard Covergroups
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

//------------ Assuming it right for time being --------------

`define RAMBASEADDR 32'h80000000
`define LARGESTPROGRAM 32'h00010000
`define SAFEREGIONSTART (`RAMBASEADDR + `LARGESTPROGRAM)
`define REGIONSTART `SAFEREGIONSTART

`define G 2              // Set G as needed (0, 1, 2, etc.)
`define g (2**(`G+2))    // Region size = 2^(G+2)

// --- STANDARD_REGION macro based on G value ---

// Case: G == 0    NA4 granularity (shift by 2)
`define REGION_G0    (`REGIONSTART >> 2)

// Case: G == 1    region has one trailing 0
`define STANDARD_REGION_G1    (`REGIONSTART >> (`G+2))

// Case: G >= 2    region has (G-1) trailing 1s
`define STANDARD_REGION_GX    (`REGIONSTART >> (`G+2)) | ((1 << (`G-1)) - 1)

// Alias one of the above depending on G
`define STANDARD_REGION `STANDARD_REGION_GX

//------------------------------------------------------------

`define COVER_RV32PMP
`define COVER_RV64PMP

covergroup PMPM_cg with function sample(ins_t ins, logic [XLEN-1:0] pmpcfg [3:0],  logic [XLEN-1:0] pmpaddr [14:0], logic [29:0] pmpcfg_rw, logic [29:0] pmpcfg_a, logic [14:0] pmpcfg_x, logic [14:0] pmpcfg_l, logic [14:0] pmp_hit);
    option.per_instance = 0;
    `include  "coverage/RISCV_coverage_standard_coverpoints.svh"

	addr_in_region: coverpoint (ins.current.rs1_val + ins.current.imm) {
    	bins at_region = {`STANDARD_REGION};
    }

    exec_instr: coverpoint ins.current.insn {
        wildcard bins jalr = {32'b????????????_?????_000_?????_1100111};
    }

    read_instr: coverpoint ins.current.insn {
        wildcard bins lb  = {32'b????????????_?????_000_?????_0000011};
        wildcard bins lbu = {32'b????????????_?????_100_?????_0000011};
        wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
        wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
        wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
        `ifdef XLEN64
            wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
            wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
        `endif
    }

    write_instr: coverpoint ins.current.insn {
        wildcard bins sb = {32'b???????_?????_?????_000_?????_0100011};
        wildcard bins sh = {32'b???????_?????_?????_001_?????_0100011};
        wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
        `ifdef XLEN64
            wildcard bins sd = {32'b???????_?????_?????_011_?????_0100011};
        `endif
    }

//-------------------------------------------------------

    standard_region: coverpoint pmpaddr[0] {
        bins standard_region = {`STANDARD_REGION};
    }

    legal_lxwr: coverpoint pmpcfg[0][7:0] {
            wildcard bins cfg_l000 = {8'b10011000};
            wildcard bins cfg_l001 = {8'b10011001};
            wildcard bins cfg_l011 = {8'b10011011};
            wildcard bins cfg_l100 = {8'b10011100};
            wildcard bins cfg_l101 = {8'b10011101};
            wildcard bins cfg_l111 = {8'b10011111};
    }

    cp_cfg_X: cross priv_mode_m, legal_lxwr, exec_instr, standard_region, addr_in_region ;
    cp_cfg_R: cross priv_mode_m, legal_lxwr, read_instr, standard_region, addr_in_region ;
    cp_cfg_W: cross priv_mode_m, legal_lxwr, write_instr, standard_region, addr_in_region ;

//-------------------------------------------------------

	X0: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x0   = {75'b??????????????0_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_x0   = {75'b?????????????0?_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_x0   = {75'b????????????0??_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_x0   = {75'b???????????0???_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_x0   = {75'b??????????0????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_x0   = {75'b?????????0?????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_x0   = {75'b????????0??????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_x0   = {75'b???????0???????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_x0   = {75'b??????0????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_x0   = {75'b?????0?????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_x0  = {75'b????0??????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_x0  = {75'b???0???????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_x0  = {75'b??0????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_x0  = {75'b?0?????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_x0  = {75'b0??????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	X1: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x1   = {75'b??????????????1_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_x1   = {75'b?????????????1?_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_x1   = {75'b????????????1??_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_x1   = {75'b???????????1???_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_x1   = {75'b??????????1????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_x1   = {75'b?????????1?????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_x1   = {75'b????????1??????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_x1   = {75'b???????1???????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_x1   = {75'b??????1????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_x1   = {75'b?????1?????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_x1  = {75'b????1??????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_x1  = {75'b???1???????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_x1  = {75'b??1????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_x1  = {75'b?1?????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_x1  = {75'b1??????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	cp_cfg_X1_all: cross priv_mode_m, exec_instr, X1, addr_in_region ;
	cp_cfg_X0_all: cross priv_mode_m, exec_instr, X0, addr_in_region ;

//-------------------------------------------------------

	RW00: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw00   = {90'b????????????????????????????00_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw00   = {90'b??????????????????????????00??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw00   = {90'b????????????????????????00????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw00   = {90'b??????????????????????00??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw00   = {90'b????????????????????00????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw00   = {90'b??????????????????00??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw00   = {90'b????????????????00????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw00   = {90'b??????????????00??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw00   = {90'b????????????00????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw00   = {90'b??????????00??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw00  = {90'b????????00????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw00  = {90'b??????00??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw00  = {90'b????00????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw00  = {90'b??00??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw00  = {90'b00????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	RW11: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 3, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????11_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????11??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????11????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????11??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????11????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????11??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????11????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????11??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw11     = {90'b????????????11????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw11     = {90'b??????????11??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw11    = {90'b????????11????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw11    = {90'b??????11??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw11    = {90'b????11????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw11    = {90'b??11??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw11    = {90'b11????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	RW10: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????01_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????01??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????01????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????01??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????01????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????01??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????01????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????01??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw11     = {90'b????????????01????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw11     = {90'b??????????01??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw11    = {90'b????????01????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw11    = {90'b??????01??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw11    = {90'b????01????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw11    = {90'b??01??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw11    = {90'b01????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	cp_cfg_Rw00_all: cross priv_mode_m, read_instr, RW00, addr_in_region ;
	cp_cfg_Rw10_all: cross priv_mode_m, read_instr, RW10, addr_in_region ;
	cp_cfg_Rw11_all: cross priv_mode_m, read_instr, RW11, addr_in_region ;
	cp_cfg_rW00_all: cross priv_mode_m, write_instr, RW00, addr_in_region ;
	cp_cfg_rW10_all: cross priv_mode_m, write_instr, RW10, addr_in_region ;
	cp_cfg_rW11_all: cross priv_mode_m, write_instr, RW11, addr_in_region ;

//-------------------------------------------------------

	RWX000: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 0 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rwx000     = {105'b????????????????????????????00_??????????????0_??????????????0_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rwx000     = {105'b??????????????????????????00??_?????????????0?_?????????????0?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rwx000     = {105'b????????????????????????00????_????????????0??_????????????0??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rwx000     = {105'b??????????????????????00??????_???????????0???_???????????0???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rwx000     = {105'b????????????????????00????????_??????????0????_??????????0????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rwx000     = {105'b??????????????????00??????????_?????????0?????_?????????0?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rwx000     = {105'b????????????????00????????????_????????0??????_????????0??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rwx000     = {105'b??????????????00??????????????_???????0???????_???????0???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rwx000     = {105'b????????????00????????????????_??????0????????_??????0????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rwx000     = {105'b??????????00??????????????????_?????0?????????_?????0?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rwx000    = {105'b????????00????????????????????_????0??????????_????0??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rwx000    = {105'b??????00??????????????????????_???0???????????_???0???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rwx000    = {105'b????00????????????????????????_??0????????????_??0????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rwx000    = {105'b??00??????????????????????????_?0?????????????_?0?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rwx000    = {105'b00????????????????????????????_0??????????????_0??????????????_11????????????????????????????_100000000000000};
	}

	cp_cfg_L_access_exec: cross priv_mode_m, exec_instr, RWX000, addr_in_region ;

	cp_cfg_L_access_read: cross priv_mode_m, read_instr, RWX000, addr_in_region ;

	cp_cfg_L_access_write: cross priv_mode_m, write_instr, RWX000, addr_in_region ;

//-------------------------------------------------------

	// Lock pmp_region_1 and check the writes on pmp_region_1 and pmp_region_0
	lock_checking: coverpoint pmpcfg_l[1] {
		bins region_locked = {1'b1};
		bins region_unlocked = {1'b0};
	}

	// Setting pmp_region_1 so incase of TOR we can check lock for pmp_region_0
	pmp_region: coverpoint pmpcfg[1][12:11] {
		bins OFF   = {2'b00};
		bins TOR   = {2'b01};
		bins NAPOT = {2'b11};
	}

	pmpcfg_xwr: coverpoint ins.prev.csr[12'h3A1][6:0] { // Region 1
		bins NAPOT_XWR = {7'b0011111};
	}

	pmpaddr: coverpoint ins.prev.csr[12'h3B1] { // Region 1
		bins four = {4};
	}

	rs1_val: coverpoint ins.prev.rs1_val { // It will try to change pmpaddr_i-1 & pmpcfg_i-1 to 00000111
		bins lockoff = {7};
	}

	write_pmp_csr: coverpoint ins.prev.insn {
		wildcard bins write_pmpaddr  = {32'b001110100001_00000_010_?????_1110011}; // Try to write value of x0 in pmpaddr[1]
		wildcard bins write_pmpcfg   = {32'b001110110001_00000_010_?????_1110011}; // Try to write value of x0 in pmpcfg[1]
		wildcard bins clear_lock_bit = {32'b001110110001_?????_011_?????_1110011}; // Try to clear pmpcfg_l[1]
	}

	write_lower_pmp_csr: coverpoint ins.prev.insn {
		wildcard bins write_pmpaddr  = {32'b001110100000_?????_010_?????_1110011}; // Try to write pmpaddr[0]
		wildcard bins write_pmpcfg   = {32'b001110110000_?????_010_?????_1110011}; // Try to write pmpcfg[0]
	}

	cp_cfg_L_modify: cross lock_checking, pmp_region, write_pmp_csr, pmpcfg_xwr, pmpaddr ;
	// If pmpcfg.A = TOR and pmpcfg.L = 1, pmpaddr_i-1 will be unchange but not pmpcfg_i-1.
	cp_cfg_L_modify_TOR: cross lock_checking, pmp_region, write_lower_pmp_csr, rs1_val, pmpcfg_xwr, pmpaddr ;

//-------------------------------------------------------

	cp_pmpaddr0_walk: coverpoint pmpaddr[0] {
		bins all_zeros = {0};
		bins all_ones = {-1};
		`ifdef XLEN32
			wildcard bins walking_ones_0  = {32'b???????????????????????????????1};
			wildcard bins walking_ones_1  = {32'b??????????????????????????????1?};
			wildcard bins walking_ones_2  = {32'b?????????????????????????????1??};
			wildcard bins walking_ones_3  = {32'b????????????????????????????1???};
			wildcard bins walking_ones_4  = {32'b???????????????????????????1????};
			wildcard bins walking_ones_5  = {32'b??????????????????????????1?????};
			wildcard bins walking_ones_6  = {32'b?????????????????????????1??????};
			wildcard bins walking_ones_7  = {32'b????????????????????????1???????};
			wildcard bins walking_ones_8  = {32'b???????????????????????1????????};
			wildcard bins walking_ones_9  = {32'b??????????????????????1?????????};
			wildcard bins walking_ones_10 = {32'b?????????????????????1??????????};
			wildcard bins walking_ones_11 = {32'b????????????????????1???????????};
			wildcard bins walking_ones_12 = {32'b???????????????????1????????????};
			wildcard bins walking_ones_13 = {32'b??????????????????1?????????????};
			wildcard bins walking_ones_14 = {32'b?????????????????1??????????????};
			wildcard bins walking_ones_15 = {32'b????????????????1???????????????};
			wildcard bins walking_ones_16 = {32'b???????????????1????????????????};
			wildcard bins walking_ones_17 = {32'b??????????????1?????????????????};
			wildcard bins walking_ones_18 = {32'b?????????????1??????????????????};
			wildcard bins walking_ones_19 = {32'b????????????1???????????????????};
			wildcard bins walking_ones_20 = {32'b???????????1????????????????????};
			wildcard bins walking_ones_21 = {32'b??????????1?????????????????????};
			wildcard bins walking_ones_22 = {32'b?????????1??????????????????????};
			wildcard bins walking_ones_23 = {32'b????????1???????????????????????};
			wildcard bins walking_ones_24 = {32'b???????1????????????????????????};
			wildcard bins walking_ones_25 = {32'b??????1?????????????????????????};
			wildcard bins walking_ones_26 = {32'b?????1??????????????????????????};
			wildcard bins walking_ones_27 = {32'b????1???????????????????????????};
			wildcard bins walking_ones_28 = {32'b???1????????????????????????????};
			wildcard bins walking_ones_29 = {32'b??1?????????????????????????????};
			wildcard bins walking_ones_30 = {32'b?1??????????????????????????????};
			wildcard bins walking_ones_31 = {32'b1???????????????????????????????};
		`endif
		`ifdef XLEN64
			wildcard bins walking_ones_0  = {54'b?????????????????????????????????????????????????????1};
			wildcard bins walking_ones_1  = {54'b????????????????????????????????????????????????????1?};
			wildcard bins walking_ones_2  = {54'b???????????????????????????????????????????????????1??};
			wildcard bins walking_ones_3  = {54'b??????????????????????????????????????????????????1???};
			wildcard bins walking_ones_4  = {54'b?????????????????????????????????????????????????1????};
			wildcard bins walking_ones_5  = {54'b????????????????????????????????????????????????1?????};
			wildcard bins walking_ones_6  = {54'b???????????????????????????????????????????????1??????};
			wildcard bins walking_ones_7  = {54'b??????????????????????????????????????????????1???????};
			wildcard bins walking_ones_8  = {54'b?????????????????????????????????????????????1????????};
			wildcard bins walking_ones_9  = {54'b????????????????????????????????????????????1?????????};
			wildcard bins walking_ones_10 = {54'b???????????????????????????????????????????1??????????};
			wildcard bins walking_ones_11 = {54'b??????????????????????????????????????????1???????????};
			wildcard bins walking_ones_12 = {54'b?????????????????????????????????????????1????????????};
			wildcard bins walking_ones_13 = {54'b????????????????????????????????????????1?????????????};
			wildcard bins walking_ones_14 = {54'b???????????????????????????????????????1??????????????};
			wildcard bins walking_ones_15 = {54'b??????????????????????????????????????1???????????????};
			wildcard bins walking_ones_16 = {54'b?????????????????????????????????????1????????????????};
			wildcard bins walking_ones_17 = {54'b????????????????????????????????????1?????????????????};
			wildcard bins walking_ones_18 = {54'b???????????????????????????????????1??????????????????};
			wildcard bins walking_ones_19 = {54'b??????????????????????????????????1???????????????????};
			wildcard bins walking_ones_20 = {54'b?????????????????????????????????1????????????????????};
			wildcard bins walking_ones_21 = {54'b????????????????????????????????1?????????????????????};
			wildcard bins walking_ones_22 = {54'b???????????????????????????????1??????????????????????};
			wildcard bins walking_ones_23 = {54'b??????????????????????????????1???????????????????????};
			wildcard bins walking_ones_24 = {54'b?????????????????????????????1????????????????????????};
			wildcard bins walking_ones_25 = {54'b????????????????????????????1?????????????????????????};
			wildcard bins walking_ones_26 = {54'b???????????????????????????1??????????????????????????};
			wildcard bins walking_ones_27 = {54'b??????????????????????????1???????????????????????????};
			wildcard bins walking_ones_28 = {54'b?????????????????????????1????????????????????????????};
			wildcard bins walking_ones_29 = {54'b????????????????????????1?????????????????????????????};
			wildcard bins walking_ones_30 = {54'b???????????????????????1??????????????????????????????};
			wildcard bins walking_ones_31 = {54'b??????????????????????1???????????????????????????????};
			wildcard bins walking_ones_32 = {54'b?????????????????????1????????????????????????????????};
			wildcard bins walking_ones_33 = {54'b????????????????????1?????????????????????????????????};
			wildcard bins walking_ones_34 = {54'b???????????????????1??????????????????????????????????};
			wildcard bins walking_ones_35 = {54'b??????????????????1???????????????????????????????????};
			wildcard bins walking_ones_36 = {54'b?????????????????1????????????????????????????????????};
			wildcard bins walking_ones_37 = {54'b????????????????1?????????????????????????????????????};
			wildcard bins walking_ones_38 = {54'b???????????????1??????????????????????????????????????};
			wildcard bins walking_ones_39 = {54'b??????????????1???????????????????????????????????????};
			wildcard bins walking_ones_40 = {54'b?????????????1????????????????????????????????????????};
			wildcard bins walking_ones_41 = {54'b????????????1?????????????????????????????????????????};
			wildcard bins walking_ones_42 = {54'b???????????1??????????????????????????????????????????};
			wildcard bins walking_ones_43 = {54'b??????????1???????????????????????????????????????????};
			wildcard bins walking_ones_44 = {54'b?????????1????????????????????????????????????????????};
			wildcard bins walking_ones_45 = {54'b????????1?????????????????????????????????????????????};
			wildcard bins walking_ones_46 = {54'b???????1??????????????????????????????????????????????};
			wildcard bins walking_ones_47 = {54'b??????1???????????????????????????????????????????????};
			wildcard bins walking_ones_48 = {54'b?????1????????????????????????????????????????????????};
			wildcard bins walking_ones_49 = {54'b????1?????????????????????????????????????????????????};
			wildcard bins walking_ones_50 = {54'b???1??????????????????????????????????????????????????};
			wildcard bins walking_ones_51 = {54'b??1???????????????????????????????????????????????????};
			wildcard bins walking_ones_52 = {54'b?1????????????????????????????????????????????????????};
			wildcard bins walking_ones_53 = {54'b1?????????????????????????????????????????????????????};
		`endif
	}

	cp_pmpcfg0_walk: coverpoint pmpcfg[0] {
		`ifdef XLEN32
			wildcard bins walking_ones_0  = {32'b???????????????????????????????1};
			wildcard bins walking_ones_1  = {32'b??????????????????????????????1?};
			wildcard bins walking_ones_2  = {32'b?????????????????????????????1??};
			wildcard bins walking_ones_3  = {32'b????????????????????????????1???};
			wildcard bins walking_ones_4  = {32'b???????????????????????????1????};
			wildcard bins walking_ones_5  = {32'b??????????????????????????1?????};
			wildcard bins walking_ones_6  = {32'b?????????????????????????1??????};
			wildcard bins walking_ones_7  = {32'b????????????????????????1???????};
			wildcard bins walking_ones_8  = {32'b???????????????????????1????????};
			wildcard bins walking_ones_9  = {32'b??????????????????????1?????????};
			wildcard bins walking_ones_10 = {32'b?????????????????????1??????????};
			wildcard bins walking_ones_11 = {32'b????????????????????1???????????};
			wildcard bins walking_ones_12 = {32'b???????????????????1????????????};
			wildcard bins walking_ones_13 = {32'b??????????????????1?????????????};
			wildcard bins walking_ones_14 = {32'b?????????????????1??????????????};
			wildcard bins walking_ones_15 = {32'b????????????????1???????????????};
			wildcard bins walking_ones_16 = {32'b???????????????1????????????????};
			wildcard bins walking_ones_17 = {32'b??????????????1?????????????????};
			wildcard bins walking_ones_18 = {32'b?????????????1??????????????????};
			wildcard bins walking_ones_19 = {32'b????????????1???????????????????};
			wildcard bins walking_ones_20 = {32'b???????????1????????????????????};
			wildcard bins walking_ones_21 = {32'b??????????1?????????????????????};
			wildcard bins walking_ones_22 = {32'b?????????1??????????????????????};
			wildcard bins walking_ones_23 = {32'b????????1???????????????????????};
			wildcard bins walking_ones_24 = {32'b???????1????????????????????????};
			wildcard bins walking_ones_25 = {32'b??????1?????????????????????????};
			wildcard bins walking_ones_26 = {32'b?????1??????????????????????????};
			wildcard bins walking_ones_27 = {32'b????1???????????????????????????};
			wildcard bins walking_ones_28 = {32'b???1????????????????????????????};
			wildcard bins walking_ones_29 = {32'b??1?????????????????????????????};
			wildcard bins walking_ones_30 = {32'b?1??????????????????????????????};
			wildcard bins walking_ones_31 = {32'b1???????????????????????????????};
		`endif
		`ifdef XLEN64
			wildcard bins walking_ones_0  = {64'b???????????????????????????????????????????????????????????????1};
			wildcard bins walking_ones_1  = {64'b??????????????????????????????????????????????????????????????1?};
			wildcard bins walking_ones_2  = {64'b?????????????????????????????????????????????????????????????1??};
			wildcard bins walking_ones_3  = {64'b????????????????????????????????????????????????????????????1???};
			wildcard bins walking_ones_4  = {64'b???????????????????????????????????????????????????????????1????};
			wildcard bins walking_ones_5  = {64'b??????????????????????????????????????????????????????????1?????};
			wildcard bins walking_ones_6  = {64'b?????????????????????????????????????????????????????????1??????};
			wildcard bins walking_ones_7  = {64'b????????????????????????????????????????????????????????1???????};
			wildcard bins walking_ones_8  = {64'b???????????????????????????????????????????????????????1????????};
			wildcard bins walking_ones_9  = {64'b??????????????????????????????????????????????????????1?????????};
			wildcard bins walking_ones_10 = {64'b?????????????????????????????????????????????????????1??????????};
			wildcard bins walking_ones_11 = {64'b????????????????????????????????????????????????????1???????????};
			wildcard bins walking_ones_12 = {64'b???????????????????????????????????????????????????1????????????};
			wildcard bins walking_ones_13 = {64'b??????????????????????????????????????????????????1?????????????};
			wildcard bins walking_ones_14 = {64'b?????????????????????????????????????????????????1??????????????};
			wildcard bins walking_ones_15 = {64'b????????????????????????????????????????????????1???????????????};
			wildcard bins walking_ones_16 = {64'b???????????????????????????????????????????????1????????????????};
			wildcard bins walking_ones_17 = {64'b??????????????????????????????????????????????1?????????????????};
			wildcard bins walking_ones_18 = {64'b?????????????????????????????????????????????1??????????????????};
			wildcard bins walking_ones_19 = {64'b????????????????????????????????????????????1???????????????????};
			wildcard bins walking_ones_20 = {64'b???????????????????????????????????????????1????????????????????};
			wildcard bins walking_ones_21 = {64'b??????????????????????????????????????????1?????????????????????};
			wildcard bins walking_ones_22 = {64'b?????????????????????????????????????????1??????????????????????};
			wildcard bins walking_ones_23 = {64'b????????????????????????????????????????1???????????????????????};
			wildcard bins walking_ones_24 = {64'b???????????????????????????????????????1????????????????????????};
			wildcard bins walking_ones_25 = {64'b??????????????????????????????????????1?????????????????????????};
			wildcard bins walking_ones_26 = {64'b?????????????????????????????????????1??????????????????????????};
			wildcard bins walking_ones_27 = {64'b????????????????????????????????????1???????????????????????????};
			wildcard bins walking_ones_28 = {64'b???????????????????????????????????1????????????????????????????};
			wildcard bins walking_ones_29 = {64'b??????????????????????????????????1?????????????????????????????};
			wildcard bins walking_ones_30 = {64'b?????????????????????????????????1??????????????????????????????};
			wildcard bins walking_ones_31 = {64'b????????????????????????????????1???????????????????????????????};
			wildcard bins walking_ones_32 = {64'b???????????????????????????????1????????????????????????????????};
			wildcard bins walking_ones_33 = {64'b??????????????????????????????1?????????????????????????????????};
			wildcard bins walking_ones_34 = {64'b?????????????????????????????1??????????????????????????????????};
			wildcard bins walking_ones_35 = {64'b????????????????????????????1???????????????????????????????????};
			wildcard bins walking_ones_36 = {64'b???????????????????????????1????????????????????????????????????};
			wildcard bins walking_ones_37 = {64'b??????????????????????????1?????????????????????????????????????};
			wildcard bins walking_ones_38 = {64'b?????????????????????????1??????????????????????????????????????};
			wildcard bins walking_ones_39 = {64'b????????????????????????1???????????????????????????????????????};
			wildcard bins walking_ones_40 = {64'b???????????????????????1????????????????????????????????????????};
			wildcard bins walking_ones_41 = {64'b??????????????????????1?????????????????????????????????????????};
			wildcard bins walking_ones_42 = {64'b?????????????????????1??????????????????????????????????????????};
			wildcard bins walking_ones_43 = {64'b????????????????????1???????????????????????????????????????????};
			wildcard bins walking_ones_44 = {64'b???????????????????1????????????????????????????????????????????};
			wildcard bins walking_ones_45 = {64'b??????????????????1?????????????????????????????????????????????};
			wildcard bins walking_ones_46 = {64'b?????????????????1??????????????????????????????????????????????};
			wildcard bins walking_ones_47 = {64'b????????????????1???????????????????????????????????????????????};
			wildcard bins walking_ones_48 = {64'b???????????????1????????????????????????????????????????????????};
			wildcard bins walking_ones_49 = {64'b??????????????1?????????????????????????????????????????????????};
			wildcard bins walking_ones_50 = {64'b?????????????1??????????????????????????????????????????????????};
			wildcard bins walking_ones_51 = {64'b????????????1???????????????????????????????????????????????????};
			wildcard bins walking_ones_52 = {64'b???????????1????????????????????????????????????????????????????};
			wildcard bins walking_ones_53 = {64'b??????????1?????????????????????????????????????????????????????};
			wildcard bins walking_ones_54 = {64'b?????????1??????????????????????????????????????????????????????};
			wildcard bins walking_ones_55 = {64'b????????1???????????????????????????????????????????????????????};
			wildcard bins walking_ones_56 = {64'b???????1????????????????????????????????????????????????????????};
			wildcard bins walking_ones_57 = {64'b??????1?????????????????????????????????????????????????????????};
			wildcard bins walking_ones_58 = {64'b?????1??????????????????????????????????????????????????????????};
			wildcard bins walking_ones_59 = {64'b????1???????????????????????????????????????????????????????????};
			wildcard bins walking_ones_60 = {64'b???1????????????????????????????????????????????????????????????};
			wildcard bins walking_ones_61 = {64'b??1?????????????????????????????????????????????????????????????};
			wildcard bins walking_ones_62 = {64'b?1??????????????????????????????????????????????????????????????};
			wildcard bins walking_ones_63 = {64'b1???????????????????????????????????????????????????????????????};
		`endif
	}

endgroup

function void pmp_sample(int hart, int issue, ins_t ins);

    logic [XLEN-1:0] pmpcfg [3:0];
    logic [XLEN-1:0] pmpaddr [14:0];
    logic [29:0] pmpcfg_rw, pmpcfg_a;
    logic [14:0] pmpcfg_x, pmpcfg_l, pmp_hit;

    for (int i = 0; i < 4; i++) begin
        pmpcfg[i] = ins.current.csr[12'h3A0 + i];
    end

    for (int j = 0; j < 15; j++) begin
        pmpaddr[j] = ins.current.csr[12'h3B0 + j];
    end

	for (int k = 0; k < 15; k++) begin
	    pmp_hit[k] = (pmpaddr[k] == `REGIONSTART);
	end

	`ifdef XLEN32
		pmpcfg_rw = {
					ins.current.csr[12'h3A3][17:16],
					ins.current.csr[12'h3A3][9:8],
					ins.current.csr[12'h3A3][1:0],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A1][25:24],
					ins.current.csr[12'h3A1][17:16],
					ins.current.csr[12'h3A1][9:8],
					ins.current.csr[12'h3A1][1:0],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_rw = {
					ins.current.csr[12'h3A2][49:48],
					ins.current.csr[12'h3A2][41:40],
					ins.current.csr[12'h3A2][33:32],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A0][57:56],
					ins.current.csr[12'h3A0][49:48],
					ins.current.csr[12'h3A0][41:40],
					ins.current.csr[12'h3A0][33:32],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_x =  {
					ins.current.csr[12'h3A3][18],
					ins.current.csr[12'h3A3][10],
					ins.current.csr[12'h3A3][2],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A1][26],
					ins.current.csr[12'h3A1][18],
					ins.current.csr[12'h3A1][10],
					ins.current.csr[12'h3A1][2],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_x =  {
					ins.current.csr[12'h3A2][50],
					ins.current.csr[12'h3A2][42],
					ins.current.csr[12'h3A2][34],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A0][58],
					ins.current.csr[12'h3A0][50],
					ins.current.csr[12'h3A0][42],
					ins.current.csr[12'h3A0][34],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_a =  {
					ins.current.csr[12'h3A3][20:19],
					ins.current.csr[12'h3A3][12:11],
					ins.current.csr[12'h3A3][4:3],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A1][28:27],
					ins.current.csr[12'h3A1][20:19],
					ins.current.csr[12'h3A1][12:11],
					ins.current.csr[12'h3A1][4:3],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_a =  {
					ins.current.csr[12'h3A2][52:51],
					ins.current.csr[12'h3A2][44:43],
					ins.current.csr[12'h3A2][36:35],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A0][60:59],
					ins.current.csr[12'h3A0][52:51],
					ins.current.csr[12'h3A0][44:43],
					ins.current.csr[12'h3A0][36:35],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_l =  {
					ins.current.csr[12'h3A3][23],
					ins.current.csr[12'h3A3][15],
					ins.current.csr[12'h3A3][7],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A1][31],
					ins.current.csr[12'h3A1][23],
					ins.current.csr[12'h3A1][15],
					ins.current.csr[12'h3A1][7],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_l =  {
					ins.current.csr[12'h3A2][55],
					ins.current.csr[12'h3A2][47],
					ins.current.csr[12'h3A2][39],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A0][63],
					ins.current.csr[12'h3A0][55],
					ins.current.csr[12'h3A0][47],
					ins.current.csr[12'h3A0][39],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif

    PMPM_cg.sample(ins, pmpcfg, pmpaddr, pmpcfg_rw, pmpcfg_a, pmpcfg_x, pmpcfg_l, pmp_hit);
endfunction
