///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fcvtmod_w_d_cg = new(); fcvtmod_w_d_cg.set_inst_name("obj_fcvtmod_w_d");
    fleq_d_cg = new(); fleq_d_cg.set_inst_name("obj_fleq_d");
    fli_d_cg = new(); fli_d_cg.set_inst_name("obj_fli_d");
    fltq_d_cg = new(); fltq_d_cg.set_inst_name("obj_fltq_d");
    fmaxm_d_cg = new(); fmaxm_d_cg.set_inst_name("obj_fmaxm_d");
    fminm_d_cg = new(); fminm_d_cg.set_inst_name("obj_fminm_d");
    fround_d_cg = new(); fround_d_cg.set_inst_name("obj_fround_d");
    froundnx_d_cg = new(); froundnx_d_cg.set_inst_name("obj_froundnx_d");
