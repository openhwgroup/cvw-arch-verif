///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

RV32CBO_PMP_exceptions_cg = new(); RV32CBO_PMP_exceptions_cg.set_inst_name("obj_RV32CBO_PMP_exceptions");