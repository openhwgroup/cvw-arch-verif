///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    czero_eqz_cg = new(); czero_eqz_cg.set_inst_name("obj_czero_eqz");
    czero_nez_cg = new(); czero_nez_cg.set_inst_name("obj_czero_nez");
