///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    div_cg = new(); div_cg.set_inst_name("obj_div");
    divu_cg = new(); divu_cg.set_inst_name("obj_divu");
    mul_cg = new(); mul_cg.set_inst_name("obj_mul");
    mulh_cg = new(); mulh_cg.set_inst_name("obj_mulh");
    mulhsu_cg = new(); mulhsu_cg.set_inst_name("obj_mulhsu");
    mulhu_cg = new(); mulhu_cg.set_inst_name("obj_mulhu");
    rem_cg = new(); rem_cg.set_inst_name("obj_rem");
    remu_cg = new(); remu_cg.set_inst_name("obj_remu");
