///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    add_uw_cg = new(); add_uw_cg.set_inst_name("obj_add_uw");
    sh1add_cg = new(); sh1add_cg.set_inst_name("obj_sh1add");
    sh1add_uw_cg = new(); sh1add_uw_cg.set_inst_name("obj_sh1add_uw");
    sh2add_cg = new(); sh2add_cg.set_inst_name("obj_sh2add");
    sh2add_uw_cg = new(); sh2add_uw_cg.set_inst_name("obj_sh2add_uw");
    sh3add_cg = new(); sh3add_cg.set_inst_name("obj_sh3add");
    sh3add_uw_cg = new(); sh3add_uw_cg.set_inst_name("obj_sh3add_uw");
    slli_uw_cg = new(); slli_uw_cg.set_inst_name("obj_slli_uw");
