///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    Ssstrict_mcsr_cg = new();         Ssstrict_mcsr_cg.set_inst_name("obj_Ssstrict_mcsr");
    Ssstrict_instr_cg = new();        Ssstrict_instr_cg.set_inst_name("obj_Ssstrict_instr");
    Ssstrict_comp_instr_cg = new();   Ssstrict_comp_instr_cg.set_inst_name("obj_Ssstrict_comp_instr");
     
