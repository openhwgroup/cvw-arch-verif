///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fleq_h_cg = new(); fleq_h_cg.set_inst_name("obj_fleq_h");
    fli_h_cg = new(); fli_h_cg.set_inst_name("obj_fli_h");
    fltq_h_cg = new(); fltq_h_cg.set_inst_name("obj_fltq_h");
    fmaxm_h_cg = new(); fmaxm_h_cg.set_inst_name("obj_fmaxm_h");
    fminm_h_cg = new(); fminm_h_cg.set_inst_name("obj_fminm_h");
    fround_h_cg = new(); fround_h_cg.set_inst_name("obj_fround_h");
    froundnx_h_cg = new(); froundnx_h_cg.set_inst_name("obj_froundnx_h");
