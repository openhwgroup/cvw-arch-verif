///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    sha256sig0_cg = new(); sha256sig0_cg.set_inst_name("obj_sha256sig0");
    sha256sig1_cg = new(); sha256sig1_cg.set_inst_name("obj_sha256sig1");
    sha256sum0_cg = new(); sha256sum0_cg.set_inst_name("obj_sha256sum0");
    sha256xum1_cg = new(); sha256xum1_cg.set_inst_name("obj_sha256xum1");
    sha512sig0_cg = new(); sha512sig0_cg.set_inst_name("obj_sha512sig0");
    sha512sig1_cg = new(); sha512sig1_cg.set_inst_name("obj_sha512sig1");
    sha512sum0_cg = new(); sha512sum0_cg.set_inst_name("obj_sha512sum0");
    sha512sum1_cg = new(); sha512sum1_cg.set_inst_name("obj_sha512sum1");
