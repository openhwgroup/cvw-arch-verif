///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    c_sext_b_cg = new(); c_sext_b_cg.set_inst_name("obj_c_sext_b");
    c_sext_h_cg = new(); c_sext_h_cg.set_inst_name("obj_c_sext_h");
    c_zext_h_cg = new(); c_zext_h_cg.set_inst_name("obj_c_zext_h");
