    `include "RV64VM_coverage.sv"
    `include "RV64VM_PMP_coverage.sv"
    `include "RV64Zicbom_coverage.sv"
    `include "RV64Zicntr_coverage.sv"
    `include "RV64Zihpm_coverage.sv"
