///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    bclr_cg = new(); bclr_cg.set_inst_name("obj_bclr");
    bclri_cg = new(); bclri_cg.set_inst_name("obj_bclri");
    bext_cg = new(); bext_cg.set_inst_name("obj_bext");
    bexti_cg = new(); bexti_cg.set_inst_name("obj_bexti");
    binv_cg = new(); binv_cg.set_inst_name("obj_binv");
    binvi_cg = new(); binvi_cg.set_inst_name("obj_binvi");
    bset_cg = new(); bset_cg.set_inst_name("obj_bset");
    bseti_cg = new(); bseti_cg.set_inst_name("obj_bseti");
