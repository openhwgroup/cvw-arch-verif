///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    amoadd_d_cg = new(); amoadd_d_cg.set_inst_name("obj_amoadd_d");
    amoadd_w_cg = new(); amoadd_w_cg.set_inst_name("obj_amoadd_w");
    amoand_d_cg = new(); amoand_d_cg.set_inst_name("obj_amoand_d");
    amoand_w_cg = new(); amoand_w_cg.set_inst_name("obj_amoand_w");
    amoaxor_d_cg = new(); amoaxor_d_cg.set_inst_name("obj_amoaxor_d");
    amoaxor_w_cg = new(); amoaxor_w_cg.set_inst_name("obj_amoaxor_w");
    amomax_d_cg = new(); amomax_d_cg.set_inst_name("obj_amomax_d");
    amomax_w_cg = new(); amomax_w_cg.set_inst_name("obj_amomax_w");
    amomaxu_d_cg = new(); amomaxu_d_cg.set_inst_name("obj_amomaxu_d");
    amomaxu_w_cg = new(); amomaxu_w_cg.set_inst_name("obj_amomaxu_w");
    amomin_d_cg = new(); amomin_d_cg.set_inst_name("obj_amomin_d");
    amomin_w_cg = new(); amomin_w_cg.set_inst_name("obj_amomin_w");
    amominu_d_cg = new(); amominu_d_cg.set_inst_name("obj_amominu_d");
    amominu_w_cg = new(); amominu_w_cg.set_inst_name("obj_amominu_w");
    amoor_d_cg = new(); amoor_d_cg.set_inst_name("obj_amoor_d");
    amoor_w_cg = new(); amoor_w_cg.set_inst_name("obj_amoor_w");
    amoswap_d_cg = new(); amoswap_d_cg.set_inst_name("obj_amoswap_d");
    amoswap_w_cg = new(); amoswap_w_cg.set_inst_name("obj_amoswap_w");
