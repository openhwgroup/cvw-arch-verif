///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    aes32dsi_cg = new(); aes32dsi_cg.set_inst_name("obj_aes32dsi");
    aes32dsmi_cg = new(); aes32dsmi_cg.set_inst_name("obj_aes32dsmi");
