///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fleq_s_cg = new(); fleq_s_cg.set_inst_name("obj_fleq_s");
    fli_s_cg = new(); fli_s_cg.set_inst_name("obj_fli_s");
    fltq_s_cg = new(); fltq_s_cg.set_inst_name("obj_fltq_s");
    fmaxm_s_cg = new(); fmaxm_s_cg.set_inst_name("obj_fmaxm_s");
    fminm_s_cg = new(); fminm_s_cg.set_inst_name("obj_fminm_s");
    fround_s_cg = new(); fround_s_cg.set_inst_name("obj_fround_s");
    froundnx_s_cg = new(); froundnx_s_cg.set_inst_name("obj_froundnx_s");
