///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    sha256sig0_cg = new(); sha256sig0_cg.set_inst_name("obj_sha256sig0");
    sha256sig1_cg = new(); sha256sig1_cg.set_inst_name("obj_sha256sig1");
    sha256sum0_cg = new(); sha256sum0_cg.set_inst_name("obj_sha256sum0");
    sha256xum1_cg = new(); sha256xum1_cg.set_inst_name("obj_sha256xum1");
    sha512sig0h_cg = new(); sha512sig0h_cg.set_inst_name("obj_sha512sig0h");
    sha512sig0l_cg = new(); sha512sig0l_cg.set_inst_name("obj_sha512sig0l");
    sha512sig1h_cg = new(); sha512sig1h_cg.set_inst_name("obj_sha512sig1h");
    sha512sig1l_cg = new(); sha512sig1l_cg.set_inst_name("obj_sha512sig1l");
    sha512sum0r_cg = new(); sha512sum0r_cg.set_inst_name("obj_sha512sum0r");
    sha512sum1r_cg = new(); sha512sum1r_cg.set_inst_name("obj_sha512sum1r");
