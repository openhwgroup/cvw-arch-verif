///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    exceptionsM_cg = new();         exceptionsM_cg.set_inst_name("obj_exceptionsM");
    exceptionsInstr_cg = new();     exceptionsInstr_cg.set_inst_name("obj_exceptionsInstr");
