///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Standard Covergroups
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_RV32PMP
`define COVER_RV64PMP

covergroup PMPM_cg with function sample(
										ins_t ins,
										logic [7:0] pmpcfg [63:0],			// Per region config registers
										logic [XLEN-1:0] pmpaddr [62:0],	// 63 unpacked pmpaddress registers
										logic [16*XLEN-1:0] pack_pmpaddr,	// 16 packed pmpaddress registers
										logic [29:0] pmpcfg_wr,				// first 15 regions RW fields
										logic [95:0] pmpcfg_WR,				// next 48 regions RW fields
										logic [29:0] pmpcfg_a,				// first 15 regions A fields
										logic [95:0] pmpcfg_A,				// next 48 regions A fields
										logic [14:0] pmpcfg_x,				// first 15 regions X fields
										logic [47:0] pmpcfg_X,				// next 48 regions X fields
										logic [14:0] pmpcfg_l,				// first 15 regions L fields
										logic [47:0] pmpcfg_L,				// next 48 regions L fields
										logic [14:0] pmp_hit,				// for first 15 regions indicating hit of pmp_entry
										logic [47:0] pmp_HIT				// for next 48 regions indicating hit of pmp_entry
										);
	option.per_instance = 0;
	`include  "coverage/RISCV_coverage_standard_coverpoints.svh"

	addr_in_region: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins at_region = {`REGIONSTART};
	}

	addr_offset_cp_cfg_A_napot_all: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins at_base      = {`REGIONSTART};
		bins below_base   = {`REGIONSTART-4};
		bins just_beyond  = {`REGIONSTART+`g};
	}

	address_offsets: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins at_base      = {`REGIONSTART};
		bins below_base   = {`REGIONSTART-4};
		bins above_base   = {`REGIONSTART+4};
		bins just_beyond  = {`REGIONSTART+`g};
		bins highest_word  = {`REGIONSTART +`g-4};
	}

	`ifdef G_IS_0
		addr_offset_cp_cfg_A_na4: coverpoint (ins.current.rs1_val + ins.current.imm) {
			bins at_base     = {`REGIONSTART};
			bins just_beyond = {`REGIONSTART+4};
			bins below_base  = {`REGIONSTART-4};
		}
	`endif

	addr_offset_cp_cfg_A_tor0: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins at_base      = {`REGIONSTART};
		bins below_base   = {`REGIONSTART-4};
	}

	exec_instr: coverpoint ins.current.insn {
		wildcard bins jalr = {32'b????????????_?????_000_?????_1100111};
	}

	read_instr_lw: coverpoint ins.current.insn {
		wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
	}

	read_instr: coverpoint ins.current.insn {
		wildcard bins lb  = {32'b????????????_?????_000_?????_0000011};
		wildcard bins lbu = {32'b????????????_?????_100_?????_0000011};
		wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
		wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
		wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
		`ifdef XLEN64
			wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
			wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
		`endif
	}

	read_instr_for_misaligned: coverpoint ins.current.insn {
		wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
		wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
		wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
		`ifdef XLEN64
			wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
			wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
		`endif
	}

	write_instr_sw: coverpoint ins.current.insn {
		wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
	}

	write_instr: coverpoint ins.current.insn {
		wildcard bins sb = {32'b???????_?????_?????_000_?????_0100011};
		wildcard bins sh = {32'b???????_?????_?????_001_?????_0100011};
		wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
		`ifdef XLEN64
			wildcard bins sd = {32'b???????_?????_?????_011_?????_0100011};
		`endif
	}

	write_instr_for_misaligned: coverpoint ins.current.insn {
		wildcard bins sh = {32'b???????_?????_?????_001_?????_0100011};
		wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
		`ifdef XLEN64
			wildcard bins sd = {32'b???????_?????_?????_011_?????_0100011};
		`endif
	}

//-------------------------------------------------------

	legal_lxwr: coverpoint {pmpcfg[0],pmpcfg[1],pmpcfg[2],pmpcfg[3],pmpcfg[4],pmpcfg[5],pmp_hit[5:0]} {
		wildcard bins cfg_l000 = {54'b????????????????????????????????????????10011000_100000};
		wildcard bins cfg_l001 = {54'b????????????????????????????????10011001????????_?10000};
		wildcard bins cfg_l011 = {54'b????????????????????????10011011????????????????_??1000};
		wildcard bins cfg_l100 = {54'b????????????????10011100????????????????????????_???100};
		wildcard bins cfg_l101 = {54'b????????10011101????????????????????????????????_????10};
		wildcard bins cfg_l111 = {54'b10011111????????????????????????????????????????_?????1};
	}

//-------------------------------------------------------
	// Addresses for TOR regions moving up by g*i
	addr_for_tor_all_region0: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {`REGIONSTART-4}; // Region with XWR-111 for test to be executed.
	}
	// Access at the start of the region
	addr_for_tor_all_region1: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART)};
	}
	addr_for_tor_all_region2: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + `g)};
	}
	addr_for_tor_all_region3: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 3*`g)};
	}
	addr_for_tor_all_region4: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 6*`g)};
	}
	addr_for_tor_all_region5: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 10*`g)};
	}
	addr_for_tor_all_region6: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 15*`g)};
	}
	addr_for_tor_all_region7: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 21*`g)};
	}
	addr_for_tor_all_region8: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 28*`g)};
	}
	addr_for_tor_all_region9: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 36*`g)};
	}
	addr_for_tor_all_region10: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 45*`g)};
	}
	addr_for_tor_all_region11: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 55*`g)};
	}
	addr_for_tor_all_region12: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 66*`g)};
	}
	addr_for_tor_all_region13: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 78*`g)};
	}
	addr_for_tor_all_region14: coverpoint(ins.current.rs1_val+ ins.current.imm){
		bins address = {(`REGIONSTART + 91*`g)};
	}

	// TOR regions increasing size by g*i
	pmpaddr_for_tor_region0: coverpoint (pmpaddr[0]==(`REGIONSTART >> 2))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region1: coverpoint ((pmpaddr[1]==((`REGIONSTART + 1*`g) >> 2)) && (pmpaddr[0]==(`REGIONSTART >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region2: coverpoint ((pmpaddr[2]==((`REGIONSTART + 3*`g) >> 2)) && (pmpaddr[1]==((`REGIONSTART + 1*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region3: coverpoint ((pmpaddr[3]==((`REGIONSTART + 6*`g) >> 2)) && (pmpaddr[2]==((`REGIONSTART + 3*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region4: coverpoint ((pmpaddr[4]==((`REGIONSTART + 10*`g) >> 2)) && (pmpaddr[3]==((`REGIONSTART + 6*`g) >> 2))) {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region5: coverpoint ((pmpaddr[5]==((`REGIONSTART + 15*`g) >> 2)) && (pmpaddr[4]==((`REGIONSTART + 10*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region6: coverpoint ((pmpaddr[6]==((`REGIONSTART + 21*`g) >> 2)) && (pmpaddr[5]==((`REGIONSTART + 15*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region7: coverpoint ((pmpaddr[7]==((`REGIONSTART + 28*`g) >> 2)) && (pmpaddr[6]==((`REGIONSTART + 21*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region8: coverpoint ((pmpaddr[8]==((`REGIONSTART + 36*`g) >> 2)) && (pmpaddr[7]==((`REGIONSTART + 28*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region9: coverpoint ((pmpaddr[9]==((`REGIONSTART + 45*`g) >> 2)) && (pmpaddr[8]==((`REGIONSTART + 36*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region10: coverpoint ((pmpaddr[10]==((`REGIONSTART + 55*`g) >> 2)) && (pmpaddr[9]==((`REGIONSTART + 45*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region11: coverpoint ((pmpaddr[11]==((`REGIONSTART + 66*`g) >> 2)) && (pmpaddr[10]==((`REGIONSTART + 55*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region12: coverpoint ((pmpaddr[12]==((`REGIONSTART + 78*`g) >> 2)) && (pmpaddr[11]==((`REGIONSTART + 66*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region13: coverpoint ((pmpaddr[13]==((`REGIONSTART + 91*`g) >> 2)) && (pmpaddr[12]==((`REGIONSTART + 78*`g) >> 2)))  {
		bins region_setup  = {1};
 	}
	pmpaddr_for_tor_region14: coverpoint ((pmpaddr[14]==((`REGIONSTART + 105*`g) >> 2)) && (pmpaddr[13]==((`REGIONSTART + 91*`g) >> 2)))  {
		bins region_setup  = {1};
 	}

   //15 configurtions, with  pmpcfg.L = 1, pmpcfg.A = TOR, pmpcfg.XWR=00(i%2)

 	// Region from 0 to REGIONSTART needs XWR Permissions for test to be exexcuted.
    RWXL_i111_pmp0cfg: coverpoint { pmpcfg[0]} {
   		bins pmp0cfg_wrx111  = {8'b10001111};
   }

	RWXL_i001_pmp1cfg: coverpoint pmpcfg[1] {
   		bins pmp1cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp2cfg: coverpoint pmpcfg[2] {
   		bins pmp2cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp3cfg: coverpoint pmpcfg[3] {
   		bins pmp3cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp4cfg: coverpoint pmpcfg[4] {
   		bins pmp4cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp5cfg: coverpoint pmpcfg[5] {
   		bins pmp5cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp6cfg: coverpoint pmpcfg[6] {
   		bins pmp6cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp7cfg: coverpoint pmpcfg[7] {
   		bins pmp7cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp8cfg: coverpoint pmpcfg[8] {
   		bins pmp8cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp9cfg: coverpoint pmpcfg[9] {
   		bins pmp9cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp10cfg: coverpoint pmpcfg[10] {
   		bins pmp10cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp11cfg: coverpoint pmpcfg[11] {
   		bins pmp11cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp12cfg: coverpoint pmpcfg[12] {
   		bins pmp0cfg_xwr000  = {8'b10001000};
   }

	RWXL_i001_pmp13cfg: coverpoint pmpcfg[13] {
   		bins pmp0cfg_xwr001  = {8'b10001001};
   }

	RWXL_i001_pmp14cfg: coverpoint pmpcfg[14] {
   		bins pmp0cfg_xwr000  = {8'b10001000};
   }

//-------------------------------------------------------

	pmpcfgA_OFF: coverpoint {pmpcfg_a,pmpcfg_l,pmpcfg_x,pmpcfg_wr,pmp_hit} {
		wildcard bins OFF0  = {105'b????????????????????????????00_??????????????1_??????????????0_????????????????????????????00_??????????????1};
		wildcard bins OFF1  = {105'b??????????????????????????00??_?????????????1?_?????????????0?_??????????????????????????00??_?????????????10};
		wildcard bins OFF2  = {105'b????????????????????????00????_????????????1??_????????????0??_????????????????????????00????_????????????100};
		wildcard bins OFF3  = {105'b??????????????????????00??????_???????????1???_???????????0???_??????????????????????00??????_???????????1000};
		wildcard bins OFF4  = {105'b????????????????????00????????_??????????1????_??????????0????_????????????????????00????????_??????????10000};
		wildcard bins OFF5  = {105'b??????????????????00??????????_?????????1?????_?????????0?????_??????????????????00??????????_?????????100000};
		wildcard bins OFF6  = {105'b????????????????00????????????_????????1??????_????????0??????_????????????????00????????????_????????1000000};
		wildcard bins OFF7  = {105'b??????????????00??????????????_???????1???????_???????0???????_??????????????00??????????????_???????10000000};
		wildcard bins OFF8  = {105'b????????????00????????????????_??????1????????_??????0????????_????????????00????????????????_??????100000000};
		wildcard bins OFF9  = {105'b??????????00??????????????????_?????1?????????_?????0?????????_??????????00??????????????????_?????1000000000};
		wildcard bins OFF10 = {105'b????????00????????????????????_????1??????????_????0??????????_????????00????????????????????_????10000000000};
		wildcard bins OFF11 = {105'b??????00??????????????????????_???1???????????_???0???????????_??????00??????????????????????_???100000000000};
		wildcard bins OFF12 = {105'b????00????????????????????????_??1????????????_??0????????????_????00????????????????????????_??1000000000000};
		wildcard bins OFF13 = {105'b??00??????????????????????????_?1?????????????_?0?????????????_??00??????????????????????????_?10000000000000};
		wildcard bins OFF14 = {105'b00????????????????????????????_1??????????????_0??????????????_00????????????????????????????_100000000000000};
	}

	`ifdef G_IS_0
		pmpcfgA_NA4: coverpoint {pmpcfg_a,pmpcfg_l,pmpcfg_x,pmpcfg_wr,pmp_hit} {
			wildcard bins NA40  = {105'b????????????????????????????10_??????????????1_??????????????0_????????????????????????????00_??????????????1};
			wildcard bins NA41  = {105'b??????????????????????????10??_?????????????1?_?????????????0?_??????????????????????????00??_?????????????10};
			wildcard bins NA42  = {105'b????????????????????????10????_????????????1??_????????????0??_????????????????????????00????_????????????100};
			wildcard bins NA43  = {105'b??????????????????????10??????_???????????1???_???????????0???_??????????????????????00??????_???????????1000};
			wildcard bins NA44  = {105'b????????????????????10????????_??????????1????_??????????0????_????????????????????00????????_??????????10000};
			wildcard bins NA45  = {105'b??????????????????10??????????_?????????1?????_?????????0?????_??????????????????00??????????_?????????100000};
			wildcard bins NA46  = {105'b????????????????10????????????_????????1??????_????????0??????_????????????????00????????????_????????1000000};
			wildcard bins NA47  = {105'b??????????????10??????????????_???????1???????_???????0???????_??????????????00??????????????_???????10000000};
			wildcard bins NA48  = {105'b????????????10????????????????_??????1????????_??????0????????_????????????00????????????????_??????100000000};
			wildcard bins NA49  = {105'b??????????10??????????????????_?????1?????????_?????0?????????_??????????00??????????????????_?????1000000000};
			wildcard bins NA410 = {105'b????????10????????????????????_????1??????????_????0??????????_????????00????????????????????_????10000000000};
			wildcard bins NA411 = {105'b??????10??????????????????????_???1???????????_???0???????????_??????00??????????????????????_???100000000000};
			wildcard bins NA412 = {105'b????10????????????????????????_??1????????????_??0????????????_????00????????????????????????_??1000000000000};
			wildcard bins NA413 = {105'b??10??????????????????????????_?1?????????????_?0?????????????_??00??????????????????????????_?10000000000000};
			wildcard bins NA414 = {105'b10????????????????????????????_1??????????????_0??????????????_00????????????????????????????_100000000000000};
		}
	`endif

	pmpcfgA_NAPOT: coverpoint {pmpcfg_a,pmpcfg_l,pmpcfg_x,pmpcfg_wr,pmp_hit} {
		wildcard bins NAPOT0  = {105'b????????????????????????????11_??????????????1_??????????????0_????????????????????????????00_??????????????1};
		wildcard bins NAPOT1  = {105'b??????????????????????????11??_?????????????1?_?????????????0?_??????????????????????????00??_?????????????10};
		wildcard bins NAPOT2  = {105'b????????????????????????11????_????????????1??_????????????0??_????????????????????????00????_????????????100};
		wildcard bins NAPOT3  = {105'b??????????????????????11??????_???????????1???_???????????0???_??????????????????????00??????_???????????1000};
		wildcard bins NAPOT4  = {105'b????????????????????11????????_??????????1????_??????????0????_????????????????????00????????_??????????10000};
		wildcard bins NAPOT5  = {105'b??????????????????11??????????_?????????1?????_?????????0?????_??????????????????00??????????_?????????100000};
		wildcard bins NAPOT6  = {105'b????????????????11????????????_????????1??????_????????0??????_????????????????00????????????_????????1000000};
		wildcard bins NAPOT7  = {105'b??????????????11??????????????_???????1???????_???????0???????_??????????????00??????????????_???????10000000};
		wildcard bins NAPOT8  = {105'b????????????11????????????????_??????1????????_??????0????????_????????????00????????????????_??????100000000};
		wildcard bins NAPOT9  = {105'b??????????11??????????????????_?????1?????????_?????0?????????_??????????00??????????????????_?????1000000000};
		wildcard bins NAPOT10 = {105'b????????11????????????????????_????1??????????_????0??????????_????????00????????????????????_????10000000000};
		wildcard bins NAPOT11 = {105'b??????11??????????????????????_???1???????????_???0???????????_??????00??????????????????????_???100000000000};
		wildcard bins NAPOT12 = {105'b????11????????????????????????_??1????????????_??0????????????_????00????????????????????????_??1000000000000};
		wildcard bins NAPOT13 = {105'b??11??????????????????????????_?1?????????????_?0?????????????_??00??????????????????????????_?10000000000000};
		wildcard bins NAPOT14 = {105'b11????????????????????????????_1??????????????_0??????????????_00????????????????????????????_100000000000000};
	}
//-------------------------------------------------------
	`ifndef G_IS_0
		pmpcfg0_A_mode_was_OFF: coverpoint {ins.prev.csr[12'h3A0]} {
  			wildcard bins OFF = {8'b00000???};
		}

		pmpcfg0_A_mode_was_NAPOT: coverpoint {ins.prev.csr[12'h3A0]} {
  			wildcard bins OFF = {8'b00011???};
		}

		pmpcfg0_A_mode_is_OFF: coverpoint {ins.current.csr[12'h3A0]} {
  			wildcard bins OFF = {8'b00000???};
		}

		pmpcfg0_A_mode_is_NAPOT: coverpoint {ins.current.csr[12'h3A0]} {
  			wildcard bins OFF = {8'b00011???};
		}

		pmpcfg0_A_mode_is_TOR: coverpoint {ins.current.csr[12'h3A0]} {
  			wildcard bins OFF = {8'b00001???};
		}
	`endif

	pmpcfg_for_cp_grain_check: coverpoint pmpcfg[0] {
		bins zero = {0};
	}

	pmpaddr0_for_cp_grain_check: coverpoint ins.prev.rs1_val {
		bins one = {{(`XLEN){1'b1}}};
	}

	csrrw_to_pmpaddr0: coverpoint ins.prev.insn {
		wildcard bins csrrw  = {32'b001110110000_?????_001_?????_1110011}; // A write is being performed to pmpaddr[0]
	}

	csrr_to_pmpaddr0: coverpoint ins.current.insn {
		wildcard bins csrr  = {32'b001110110000_00000_010_?????_1110011}; // A read is being performed to pmpaddr[0]
	}

//-------------------------------------------------------

	pmpcfg_for_tor0: coverpoint {pmpcfg[0]} {
		wildcard bins pmp0cfg_xwr000  = {8'b10001111}; //L=1,A=TOR,XWR=111
	}

	pmpcfg_tor_bot_L0: coverpoint ({pmpcfg[1],pmpcfg[0]}) {
    	bins pmp_cfg_tor1 =  {16'b10001101_00000000}; //L=0 for pmpcfg0 and L=1 for pmpcfg1.A=TOR,XWR=101 and 000 respectively
	}

	pmpcfg_tor_bot_L1: coverpoint ({pmpcfg[1],pmpcfg[0]}) {
		bins pmp_cfg_tor1 =  {16'b10001101_10000000}; //L=1 for pmpcfg0 and L=1 for pmpcfg1.A=TOR,XWR=101 and 000 respectively
	}

	pmp_addr_for_tor: coverpoint {pmpaddr[1],pmpaddr[0]} {
		bins range = {`NON_STANDARD_REGION+`g,`NON_STANDARD_REGION};
	}

	pmp_addr_for_tor_bot: coverpoint ({pmpaddr[1],pmpaddr[0]} == {(`REGIONSTART+`g)>>2,`REGIONSTART>>2})  {  //pmpaddr0 = pmpaddr1-g
		bins range = {1};
	}

	pmp_addr_for_tor0: coverpoint {pmpaddr[0]} {
		bins range = {`NON_STANDARD_REGION};
	}

	addr_for_tor_bot: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins pmpaddr0_4 = {((`NON_STANDARD_REGION)<<2)-4}; //pmpaddr0-4
		bins pmpaddr0 = {(`NON_STANDARD_REGION)<<2}; //pmpaddr0
		bins pmpaddr1_4 = {(`REGIONSTART+`g)-4}; //pmpaddr1-4 NOTE: REGIONSTART>>2 => NON_STANDARD_REGION (pmp encoded address)
		bins pmpaddr1 = {`REGIONSTART+`g};
	}

	pmp_addr_for_tor_nonoverlap1: coverpoint ({pmpaddr[1], pmpaddr[0]}=={`REGIONSTART>>2, `REGIONSTART>>2}) { // pmpaddr0 >= pmpaddr1.
  		bins range1 = {1};
 	}

	pmp_addr_for_tor_nonoverlap2: coverpoint ({pmpaddr[1], pmpaddr[0]}=={`REGIONSTART>>2, (`REGIONSTART+`g)>>2}) { // pmpaddr0 >= pmpaddr1.
		bins range2 = {1};
 	}

	pmp_addr_for_tor_nonoverlap3: coverpoint ({pmpaddr[1], pmpaddr[0]}=={`REGIONSTART>>2, {$bits(pmpaddr[0]){1'b1}}}) { // pmpaddr0 >= pmpaddr1.
		bins range3 = {1}; //pmpaddr0 = all 1s
 	}

	pmpcfg_tor_nonoverlap: coverpoint {pmpcfg[1],pmpcfg[0]} {
    	bins pmp_cfg_tor1 =  {16'b10001000_00000000}; //L=1 for pmpcfg1 and L=0 for pmpcfg0,A=TOR for cf1 and A=OFF for 0,XWR=000(both)
	}

	addr_for_tor_nonoverlap: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins addr1 = {(`NON_STANDARD_REGION)<<2}; //pmpaddr1
		bins addr2 = {((`NON_STANDARD_REGION)<<2)+4}; //pmpaddr1+4
		bins addr3 = {((`NON_STANDARD_REGION)<<2)-4}; //pmpaddr1-4
	}

	pmpaddr_for_napot_misaligned: coverpoint {pmpaddr[0]} {
		bins pmpaddr = {(`REGIONSTART>>2) | ((1 << (`k)) - 1) }; //No of Trailing 1s = (1 << G-1) - 1, a standard NAPOT Region
	}

	pmpcfg_for_napot_misaligned: coverpoint {pmpcfg[0]} {
		bins pmp_cfg_napot_locked = {8'b10011111}; //L=1,A=NAPOT,XWR=111
		bins pmp_cfg_napot_unlocked = {8'b00011111}; //L=0,A=NAPOT,XWR=111
	}

	pmpaddr_for_na4_misaligned: coverpoint {pmpaddr[0]} {
		bins pmpaddr = {`NON_STANDARD_REGION};
	}

	pmpcfg_for_na4_misaligned: coverpoint {pmpcfg[0]} {
		bins pmp_cfg_na4_locked = {8'b10010111}; //L=1,A=NA4,XWR=111
		bins pmp_cfg_na4_unlocked = {8'b00010111}; //L=0,A=NA4,XWR=111
	}

	addr_for_na4_misaligned_straddling_start: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins addr1 = {`REGIONSTART-1}; //for 1 byte outside the region
	}

	addr_for_na4_misaligned_straddling_end: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins addr1 = {`REGIONSTART+3}; //for 3 byte outside the region
	}

	pmpaddr_for_tor_misaligned: coverpoint ({pmpaddr[3],pmpaddr[2]}=={(`REGIONSTART+`g)>>2,`REGIONSTART>>2}) {
		bins pmpaddr = {1};
	}

	pmpcfg_for_tor_misaligned: coverpoint {pmpcfg[3]} {
		bins pmp_cfg_tor_locked = {8'b10001111}; //L=1,A=TOR,XWR=111
		bins pmp_cfg_tor_unlocked = {8'b00001111}; //L=0,A=TOR,XWR=111
	}

	addr_for_misaligned_straddling_start: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins addr1 = {`REGIONSTART-1};
	}

	addr_for_misaligned_straddling_end: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins addr1 = {(`REGIONSTART+`g)-1};
	}

	pmpcfg_for_off_misaligned: coverpoint {ins.current.csr[12'h3A0][7:0]} {
		bins pmp_cfg_tor_locked = {8'b10000111}; //L=1,A=OFF,XWR=111
		bins pmp_cfg_tor_unlocked = {8'b00000111}; //L=0,A=OFF,XWR=111
	}

	pmpaddr_for_off_misaligned: coverpoint (pmpaddr[0]==`REGIONSTART>>2) {
		bins pmpaddr = {1};
	}

//-------------------------------------------------------

	//6 legal combinations for XRW

	// Configuration for pairs of pmpaddr ((11,10),(9,8),(7,6),(5,4),(3,2),(1,0)) for Default TOR.
  	legal_RWX_L_TOR: coverpoint {pmpcfg_l[11:0], pmpcfg_a[23:0], pmpcfg_x[11:0], pmpcfg_wr[23:0], pmp_hit[11:0]} { // pmpcfg.RWX = legal combinations, pmpcfg.L = 1 and pmpcfg.A = 1
		wildcard bins pmp1cfg_lxwr_1000  = {84'b1???????????_01??????????????????????_0???????????_00??????????????????????_?1??????????};
		wildcard bins pmp1cfg_lxwr_1001  = {84'b??1?????????_????01??????????????????_??0?????????_????01??????????????????_???1????????};
		wildcard bins pmp0cfg_lxwr_1011  = {84'b????1???????_????????01??????????????_????0???????_????????11??????????????_?????1??????};
		wildcard bins pmp0cfg_lxwr_1100  = {84'b??????1?????_????????????01??????????_??????1?????_????????????00??????????_???????1????};
		wildcard bins pmp0cfg_lxwr_1101  = {84'b????????1???_????????????????01??????_????????1???_????????????????01??????_?????????1??};
		wildcard bins pmp0cfg_lxwr_1111  = {84'b??????????1?_????????????????????01??_??????????1?_????????????????????11??_???????????1};
	}

  	legal_RWX_L_NAPOT: coverpoint {pmpcfg_l[5:0], pmpcfg_a[11:0], pmpcfg_x[5:0], pmpcfg_wr[11:0], pmp_hit[5:0]} { // pmpcfg.RWX = legal combinations, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp1cfg_lxwr_1000  = {42'b1?????_11??????????_0?????_00??????????_100000};
		wildcard bins pmp1cfg_lxwr_1001  = {42'b?1????_??11????????_?0????_??01????????_?10000};
		wildcard bins pmp0cfg_lxwr_1011  = {42'b??1???_????11??????_??0???_????11??????_??1000};
		wildcard bins pmp0cfg_lxwr_1100  = {42'b???1??_??????11????_???1??_??????00????_???100};
		wildcard bins pmp0cfg_lxwr_1101  = {42'b????1?_????????11??_????1?_????????01??_????10};
		wildcard bins pmp0cfg_lxwr_1111  = {42'b?????1_??????????11_?????1_??????????11_?????1};
	}

//-------------------------------------------------------

	`ifdef G_IS_0
  		legal_RWX_L_NA4: coverpoint {pmpcfg_l[5:0], pmpcfg_a[11:0], pmpcfg_x[5:0], pmpcfg_wr[11:0], pmp_hit[5:0]} { // pmpcfg.RWX = legal combinations, pmpcfg.L = 1 and pmpcfg.A = 2'b10
			wildcard bins pmp1cfg_lxwr_1000  = {42'b1?????_10??????????_0?????_00??????????_100000};
			wildcard bins pmp1cfg_lxwr_1001  = {42'b?1????_??10????????_?0????_??01????????_?10000};
			wildcard bins pmp0cfg_lxwr_1011  = {42'b??1???_????10??????_??0???_????11??????_??1000};
			wildcard bins pmp0cfg_lxwr_1100  = {42'b???1??_??????10????_???1??_??????00????_???100};
			wildcard bins pmp0cfg_lxwr_1101  = {42'b????1?_????????10??_????1?_????????01??_????10};
			wildcard bins pmp0cfg_lxwr_1111  = {42'b?????1_??????????10_?????1_??????????11_?????1};
		}
	`endif

//-------------------------------------------------------

	X0: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x0   = {75'b??????????????0_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_x0   = {75'b?????????????0?_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_x0   = {75'b????????????0??_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_x0   = {75'b???????????0???_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_x0   = {75'b??????????0????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_x0   = {75'b?????????0?????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_x0   = {75'b????????0??????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_x0   = {75'b???????0???????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_x0   = {75'b??????0????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_x0   = {75'b?????0?????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_x0  = {75'b????0??????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_x0  = {75'b???0???????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_x0  = {75'b??0????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_x0  = {75'b?0?????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_x0  = {75'b0??????????????_1??????????????_11????????????????????????????_1??????????????};
	}

	X1: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x1   = {75'b??????????????1_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_x1   = {75'b?????????????1?_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_x1   = {75'b????????????1??_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_x1   = {75'b???????????1???_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_x1   = {75'b??????????1????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_x1   = {75'b?????????1?????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_x1   = {75'b????????1??????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_x1   = {75'b???????1???????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_x1   = {75'b??????1????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_x1   = {75'b?????1?????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_x1  = {75'b????1??????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_x1  = {75'b???1???????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_x1  = {75'b??1????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_x1  = {75'b?1?????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_x1  = {75'b1??????????????_1??????????????_11????????????????????????????_1??????????????};
	}

//-------------------------------------------------------

	RW00: coverpoint {pmpcfg_wr, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw00   = {90'b????????????????????????????00_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw00   = {90'b??????????????????????????00??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw00   = {90'b????????????????????????00????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw00   = {90'b??????????????????????00??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw00   = {90'b????????????????????00????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw00   = {90'b??????????????????00??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw00   = {90'b????????????????00????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw00   = {90'b??????????????00??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw00   = {90'b????????????00????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw00   = {90'b??????????00??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw00  = {90'b????????00????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw00  = {90'b??????00??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw00  = {90'b????00????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw00  = {90'b??00??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw00  = {90'b00????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}

	RW11: coverpoint {pmpcfg_wr, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 3, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????11_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????11??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????11????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????11??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????11????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????11??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????11????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????11??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw11     = {90'b????????????11????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw11     = {90'b??????????11??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw11    = {90'b????????11????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw11    = {90'b??????11??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw11    = {90'b????11????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw11    = {90'b??11??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw11    = {90'b11????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}

	RW10: coverpoint {pmpcfg_wr, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw10     = {90'b????????????????????????????01_??????????????1_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rw10     = {90'b??????????????????????????01??_?????????????1?_??????????????????????????11??_?????????????1?};
		wildcard bins pmp2cfg_rw10     = {90'b????????????????????????01????_????????????1??_????????????????????????11????_????????????1??};
		wildcard bins pmp3cfg_rw10     = {90'b??????????????????????01??????_???????????1???_??????????????????????11??????_???????????1???};
		wildcard bins pmp4cfg_rw10     = {90'b????????????????????01????????_??????????1????_????????????????????11????????_??????????1????};
		wildcard bins pmp5cfg_rw10     = {90'b??????????????????01??????????_?????????1?????_??????????????????11??????????_?????????1?????};
		wildcard bins pmp6cfg_rw10     = {90'b????????????????01????????????_????????1??????_????????????????11????????????_????????1??????};
		wildcard bins pmp7cfg_rw10     = {90'b??????????????01??????????????_???????1???????_??????????????11??????????????_???????1???????};
		wildcard bins pmp8cfg_rw10     = {90'b????????????01????????????????_??????1????????_????????????11????????????????_??????1????????};
		wildcard bins pmp9cfg_rw10     = {90'b??????????01??????????????????_?????1?????????_??????????11??????????????????_?????1?????????};
		wildcard bins pmp10cfg_rw10    = {90'b????????01????????????????????_????1??????????_????????11????????????????????_????1??????????};
		wildcard bins pmp11cfg_rw10    = {90'b??????01??????????????????????_???1???????????_??????11??????????????????????_???1???????????};
		wildcard bins pmp12cfg_rw10    = {90'b????01????????????????????????_??1????????????_????11????????????????????????_??1????????????};
		wildcard bins pmp13cfg_rw10    = {90'b??01??????????????????????????_?1?????????????_??11??????????????????????????_?1?????????????};
		wildcard bins pmp14cfg_rw10    = {90'b01????????????????????????????_1??????????????_11????????????????????????????_1??????????????};
	}

//-------------------------------------------------------

	RWX000: coverpoint {pmpcfg_wr, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 0 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rwx000  = {105'b????????????????????????????00_??????????????0_??????????????0_????????????????????????????11_??????????????1};
		wildcard bins pmp1cfg_rwx000  = {105'b??????????????????????????00??_?????????????0?_?????????????0?_??????????????????????????11??_?????????????10};
		wildcard bins pmp2cfg_rwx000  = {105'b????????????????????????00????_????????????0??_????????????0??_????????????????????????11????_????????????100};
		wildcard bins pmp3cfg_rwx000  = {105'b??????????????????????00??????_???????????0???_???????????0???_??????????????????????11??????_???????????1000};
		wildcard bins pmp4cfg_rwx000  = {105'b????????????????????00????????_??????????0????_??????????0????_????????????????????11????????_??????????10000};
		wildcard bins pmp5cfg_rwx000  = {105'b??????????????????00??????????_?????????0?????_?????????0?????_??????????????????11??????????_?????????100000};
		wildcard bins pmp6cfg_rwx000  = {105'b????????????????00????????????_????????0??????_????????0??????_????????????????11????????????_????????1000000};
		wildcard bins pmp7cfg_rwx000  = {105'b??????????????00??????????????_???????0???????_???????0???????_??????????????11??????????????_???????10000000};
		wildcard bins pmp8cfg_rwx000  = {105'b????????????00????????????????_??????0????????_??????0????????_????????????11????????????????_??????100000000};
		wildcard bins pmp9cfg_rwx000  = {105'b??????????00??????????????????_?????0?????????_?????0?????????_??????????11??????????????????_?????1000000000};
		wildcard bins pmp10cfg_rwx000 = {105'b????????00????????????????????_????0??????????_????0??????????_????????11????????????????????_????10000000000};
		wildcard bins pmp11cfg_rwx000 = {105'b??????00??????????????????????_???0???????????_???0???????????_??????11??????????????????????_???100000000000};
		wildcard bins pmp12cfg_rwx000 = {105'b????00????????????????????????_??0????????????_??0????????????_????11????????????????????????_??1000000000000};
		wildcard bins pmp13cfg_rwx000 = {105'b??00??????????????????????????_?0?????????????_?0?????????????_??11??????????????????????????_?10000000000000};
		wildcard bins pmp14cfg_rwx000 = {105'b00????????????????????????????_0??????????????_0??????????????_11????????????????????????????_100000000000000};
	}

//-------------------------------------------------------

	/* These coverpoints are for cp_cfg_L_modify & cp_cfg_L_modify_TOR and it will just tell
	 we're trying to write values in PMP CSRs when L = {0/1}, A = {OFF,TOR,NAPOT} and
	 we need to check from tests and logs that pmpcfg and pmpaddr are unwritable when
	 L = 1, and write to pmpaddr of previous region in case of TOR is also ignored.*/

	pmp_region: coverpoint ins.prev.csr[12'h3A0][12:11] {
		bins OFF   = {0};
		bins TOR   = {1};
		bins NAPOT = {3};
	}

	// L = {0/1} pmp_region_1 and check the writes on pmp_region_1 and pmp_region_0
	lock_checking: coverpoint ins.prev.csr[12'h3A0][15] {
		bins locked_region = {1};
		bins unlocked_region = {0};
	}

	// Attempt to write values in given PMP CSRs when A = {OFF/TOR/NAPOT} and L = {0/1}
	// rs1 should be x0 while writing to pmpaddr1 & pmp1cfg0 in order to write all 0s.
	// rs1 should be x4 with the value -1 which we try to write in lower pmpaddr.
	// rs1 should be x5 having 3'b111 for XWR at LSB to write in lower pmpcfg.
	pmp_csr_to_write: coverpoint ins.current.insn {
		wildcard bins pmpaddr1 = {32'b001110110001_00000_001_?????_1110011};
		wildcard bins pmp1cfg0 = {32'b001110100000_00000_001_?????_1110011};
		wildcard bins pmp0cfg0 = {32'b001110100000_00101_001_?????_1110011};
		wildcard bins pmpaddr0 = {32'b001110110000_00100_001_?????_1110011};
	}

//-------------------------------------------------------

	cp_walk_rs1: coverpoint ins.current.rs1_val {
		`ifdef XLEN32
			wildcard bins walking_ones_0  = {32'b00000000000000000000000000000001};
			wildcard bins walking_ones_1  = {32'b00000000000000000000000000000010};
			wildcard bins walking_ones_2  = {32'b00000000000000000000000000000100};
			wildcard bins walking_ones_3  = {32'b00000000000000000000000000001000};
			wildcard bins walking_ones_4  = {32'b00000000000000000000000000010000};
			wildcard bins walking_ones_5  = {32'b00000000000000000000000000100000};
			wildcard bins walking_ones_6  = {32'b00000000000000000000000001000000};
			wildcard bins walking_ones_7  = {32'b00000000000000000000000010000000};
			wildcard bins walking_ones_8  = {32'b00000000000000000000000100000000};
			wildcard bins walking_ones_9  = {32'b00000000000000000000001000000000};
			wildcard bins walking_ones_10 = {32'b00000000000000000000010000000000};
			wildcard bins walking_ones_11 = {32'b00000000000000000000100000000000};
			wildcard bins walking_ones_12 = {32'b00000000000000000001000000000000};
			wildcard bins walking_ones_13 = {32'b00000000000000000010000000000000};
			wildcard bins walking_ones_14 = {32'b00000000000000000100000000000000};
			wildcard bins walking_ones_15 = {32'b00000000000000001000000000000000};
			wildcard bins walking_ones_16 = {32'b00000000000000010000000000000000};
			wildcard bins walking_ones_17 = {32'b00000000000000100000000000000000};
			wildcard bins walking_ones_18 = {32'b00000000000001000000000000000000};
			wildcard bins walking_ones_19 = {32'b00000000000010000000000000000000};
			wildcard bins walking_ones_20 = {32'b00000000000100000000000000000000};
			wildcard bins walking_ones_21 = {32'b00000000001000000000000000000000};
			wildcard bins walking_ones_22 = {32'b00000000010000000000000000000000};
			wildcard bins walking_ones_23 = {32'b00000000100000000000000000000000};
			wildcard bins walking_ones_24 = {32'b00000001000000000000000000000000};
			wildcard bins walking_ones_25 = {32'b00000010000000000000000000000000};
			wildcard bins walking_ones_26 = {32'b00000100000000000000000000000000};
			wildcard bins walking_ones_27 = {32'b00001000000000000000000000000000};
			wildcard bins walking_ones_28 = {32'b00010000000000000000000000000000};
			wildcard bins walking_ones_29 = {32'b00100000000000000000000000000000};
			wildcard bins walking_ones_30 = {32'b01000000000000000000000000000000};
			wildcard bins walking_ones_31 = {32'b10000000000000000000000000000000};
		`endif
		`ifdef XLEN64
			wildcard bins walking_ones_0  = {64'b0000000000000000000000000000000000000000000000000000000000000001};
			wildcard bins walking_ones_1  = {64'b0000000000000000000000000000000000000000000000000000000000000010};
			wildcard bins walking_ones_2  = {64'b0000000000000000000000000000000000000000000000000000000000000100};
			wildcard bins walking_ones_3  = {64'b0000000000000000000000000000000000000000000000000000000000001000};
			wildcard bins walking_ones_4  = {64'b0000000000000000000000000000000000000000000000000000000000010000};
			wildcard bins walking_ones_5  = {64'b0000000000000000000000000000000000000000000000000000000000100000};
			wildcard bins walking_ones_6  = {64'b0000000000000000000000000000000000000000000000000000000001000000};
			wildcard bins walking_ones_7  = {64'b0000000000000000000000000000000000000000000000000000000010000000};
			wildcard bins walking_ones_8  = {64'b0000000000000000000000000000000000000000000000000000000100000000};
			wildcard bins walking_ones_9  = {64'b0000000000000000000000000000000000000000000000000000001000000000};
			wildcard bins walking_ones_10 = {64'b0000000000000000000000000000000000000000000000000000010000000000};
			wildcard bins walking_ones_11 = {64'b0000000000000000000000000000000000000000000000000000100000000000};
			wildcard bins walking_ones_12 = {64'b0000000000000000000000000000000000000000000000000001000000000000};
			wildcard bins walking_ones_13 = {64'b0000000000000000000000000000000000000000000000000010000000000000};
			wildcard bins walking_ones_14 = {64'b0000000000000000000000000000000000000000000000000100000000000000};
			wildcard bins walking_ones_15 = {64'b0000000000000000000000000000000000000000000000001000000000000000};
			wildcard bins walking_ones_16 = {64'b0000000000000000000000000000000000000000000000010000000000000000};
			wildcard bins walking_ones_17 = {64'b0000000000000000000000000000000000000000000000100000000000000000};
			wildcard bins walking_ones_18 = {64'b0000000000000000000000000000000000000000000001000000000000000000};
			wildcard bins walking_ones_19 = {64'b0000000000000000000000000000000000000000000010000000000000000000};
			wildcard bins walking_ones_20 = {64'b0000000000000000000000000000000000000000000100000000000000000000};
			wildcard bins walking_ones_21 = {64'b0000000000000000000000000000000000000000001000000000000000000000};
			wildcard bins walking_ones_22 = {64'b0000000000000000000000000000000000000000010000000000000000000000};
			wildcard bins walking_ones_23 = {64'b0000000000000000000000000000000000000000100000000000000000000000};
			wildcard bins walking_ones_24 = {64'b0000000000000000000000000000000000000001000000000000000000000000};
			wildcard bins walking_ones_25 = {64'b0000000000000000000000000000000000000010000000000000000000000000};
			wildcard bins walking_ones_26 = {64'b0000000000000000000000000000000000000100000000000000000000000000};
			wildcard bins walking_ones_27 = {64'b0000000000000000000000000000000000001000000000000000000000000000};
			wildcard bins walking_ones_28 = {64'b0000000000000000000000000000000000010000000000000000000000000000};
			wildcard bins walking_ones_29 = {64'b0000000000000000000000000000000000100000000000000000000000000000};
			wildcard bins walking_ones_30 = {64'b0000000000000000000000000000000001000000000000000000000000000000};
			wildcard bins walking_ones_31 = {64'b0000000000000000000000000000000010000000000000000000000000000000};
			wildcard bins walking_ones_32 = {64'b0000000000000000000000000000000100000000000000000000000000000000};
			wildcard bins walking_ones_33 = {64'b0000000000000000000000000000001000000000000000000000000000000000};
			wildcard bins walking_ones_34 = {64'b0000000000000000000000000000010000000000000000000000000000000000};
			wildcard bins walking_ones_35 = {64'b0000000000000000000000000000100000000000000000000000000000000000};
			wildcard bins walking_ones_36 = {64'b0000000000000000000000000001000000000000000000000000000000000000};
			wildcard bins walking_ones_37 = {64'b0000000000000000000000000010000000000000000000000000000000000000};
			wildcard bins walking_ones_38 = {64'b0000000000000000000000000100000000000000000000000000000000000000};
			wildcard bins walking_ones_39 = {64'b0000000000000000000000001000000000000000000000000000000000000000};
			wildcard bins walking_ones_40 = {64'b0000000000000000000000010000000000000000000000000000000000000000};
			wildcard bins walking_ones_41 = {64'b0000000000000000000000100000000000000000000000000000000000000000};
			wildcard bins walking_ones_42 = {64'b0000000000000000000001000000000000000000000000000000000000000000};
			wildcard bins walking_ones_43 = {64'b0000000000000000000010000000000000000000000000000000000000000000};
			wildcard bins walking_ones_44 = {64'b0000000000000000000100000000000000000000000000000000000000000000};
			wildcard bins walking_ones_45 = {64'b0000000000000000001000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_46 = {64'b0000000000000000010000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_47 = {64'b0000000000000000100000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_48 = {64'b0000000000000001000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_49 = {64'b0000000000000010000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_50 = {64'b0000000000000100000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_51 = {64'b0000000000001000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_52 = {64'b0000000000010000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_53 = {64'b0000000000100000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_54 = {64'b0000000001000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_55 = {64'b0000000010000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_56 = {64'b0000000100000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_57 = {64'b0000001000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_58 = {64'b0000010000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_59 = {64'b0000100000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_60 = {64'b0001000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_61 = {64'b0010000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_62 = {64'b0100000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_63 = {64'b1000000000000000000000000000000000000000000000000000000000000000};
		`endif
	}

	cp_zero_rs1: coverpoint ins.current.rs1_val {
		bins rs1_val = {0};
	}

	csrrw: coverpoint ins.current.insn {
		wildcard bins csrrw  = {32'b????????????_?????_001_?????_1110011}; // Try to write pmpaddr or pmpcfg
	}

	legal_pmpaddr_entries: coverpoint ins.current.insn[31:20] {
		bins pmpaddr0   = {12'h3B0};
		bins pmpaddr1   = {12'h3B1};
		bins pmpaddr2   = {12'h3B2};
		bins pmpaddr3   = {12'h3B3};
		bins pmpaddr4   = {12'h3B4};
		bins pmpaddr5   = {12'h3B5};
		bins pmpaddr6   = {12'h3B6};
		bins pmpaddr7   = {12'h3B7};
		bins pmpaddr8   = {12'h3B8};
		bins pmpaddr9   = {12'h3B9};
		bins pmpaddr10  = {12'h3BA};
		bins pmpaddr11  = {12'h3BB};
		bins pmpaddr12  = {12'h3BC};
		bins pmpaddr13  = {12'h3BD};
		bins pmpaddr14  = {12'h3BE};
		bins pmpaddr15  = {12'h3BF};
		`ifdef PMP_64
			bins pmpaddr16  = {12'h3C0};
			bins pmpaddr17  = {12'h3C1};
			bins pmpaddr18  = {12'h3C2};
			bins pmpaddr19  = {12'h3C3};
			bins pmpaddr20  = {12'h3C4};
			bins pmpaddr21  = {12'h3C5};
			bins pmpaddr22  = {12'h3C6};
			bins pmpaddr23  = {12'h3C7};
			bins pmpaddr24  = {12'h3C8};
			bins pmpaddr25  = {12'h3C9};
			bins pmpaddr26  = {12'h3CA};
			bins pmpaddr27  = {12'h3CB};
			bins pmpaddr28  = {12'h3CC};
			bins pmpaddr29  = {12'h3CD};
			bins pmpaddr30  = {12'h3CE};
			bins pmpaddr31  = {12'h3CF};
			bins pmpaddr32  = {12'h3D0};
			bins pmpaddr33  = {12'h3D1};
			bins pmpaddr34  = {12'h3D2};
			bins pmpaddr35  = {12'h3D3};
			bins pmpaddr36  = {12'h3D4};
			bins pmpaddr37  = {12'h3D5};
			bins pmpaddr38  = {12'h3D6};
			bins pmpaddr39  = {12'h3D7};
			bins pmpaddr40  = {12'h3D8};
			bins pmpaddr41  = {12'h3D9};
			bins pmpaddr42  = {12'h3DA};
			bins pmpaddr43  = {12'h3DB};
			bins pmpaddr44  = {12'h3DC};
			bins pmpaddr45  = {12'h3DD};
			bins pmpaddr46  = {12'h3DE};
			bins pmpaddr47  = {12'h3DF};
			bins pmpaddr48  = {12'h3E0};
			bins pmpaddr49  = {12'h3E1};
			bins pmpaddr50  = {12'h3E2};
			bins pmpaddr51  = {12'h3E3};
			bins pmpaddr52  = {12'h3E4};
			bins pmpaddr53  = {12'h3E5};
			bins pmpaddr54  = {12'h3E6};
			bins pmpaddr55  = {12'h3E7};
			bins pmpaddr56  = {12'h3E8};
			bins pmpaddr57  = {12'h3E9};
			bins pmpaddr58  = {12'h3EA};
			bins pmpaddr59  = {12'h3EB};
			bins pmpaddr60  = {12'h3EC};
			bins pmpaddr61  = {12'h3ED};
			bins pmpaddr62  = {12'h3EE};
			bins pmpaddr63  = {12'h3EF};
		`endif
	}

	legal_pmpcfg_entries_even: coverpoint ins.current.insn[31:20] { 	// For writing walking ones in even PMPCFGs
		bins pmpcfg0   = {12'h3A0};
		bins pmpcfg2   = {12'h3A2};
		`ifdef PMP_64
			bins pmpcfg4   = {12'h3A4};
			bins pmpcfg6   = {12'h3A6};
			bins pmpcfg8   = {12'h3A8};
			bins pmpcfg10  = {12'h3AA};
			bins pmpcfg12  = {12'h3AC};
			bins pmpcfg14  = {12'h3AE};
		`endif
	}

	legal_pmpcfg_entries_odd: coverpoint ins.current.insn[31:20] { 	// For writing zero in odd PMPCFGs
		bins pmpcfg1   = {12'h3A1};
		bins pmpcfg3   = {12'h3A3};
		`ifdef PMP_64
			bins pmpcfg5   = {12'h3A5};
			bins pmpcfg7   = {12'h3A7};
			bins pmpcfg9   = {12'h3A9};
			bins pmpcfg11  = {12'h3AB};
			bins pmpcfg13  = {12'h3AD};
			bins pmpcfg15  = {12'h3AF};
		`endif
	}
//-------------------------------------------------------

	`ifdef PMP_64
		pmp64: coverpoint {pmpcfg_L, pmpcfg_X, pmpcfg_wr, pmp_HIT} {
			wildcard bins pmp15cfg = {240'b???????????????????????????????????????????????1_???????????????????????????????????????????????1_??????????????????????????????????????????????????????????????????????????????????????????????01_000000000000000000000000000000000000000000000001};
			wildcard bins pmp16cfg = {240'b??????????????????????????????????????????????1?_??????????????????????????????????????????????1?_????????????????????????????????????????????????????????????????????????????????????????????01??_000000000000000000000000000000000000000000000010};
			wildcard bins pmp17cfg = {240'b?????????????????????????????????????????????1??_?????????????????????????????????????????????1??_??????????????????????????????????????????????????????????????????????????????????????????01????_000000000000000000000000000000000000000000000100};
			wildcard bins pmp18cfg = {240'b????????????????????????????????????????????1???_????????????????????????????????????????????1???_????????????????????????????????????????????????????????????????????????????????????????01??????_000000000000000000000000000000000000000000001000};
			wildcard bins pmp19cfg = {240'b???????????????????????????????????????????1????_???????????????????????????????????????????1????_??????????????????????????????????????????????????????????????????????????????????????01????????_000000000000000000000000000000000000000000010000};
			wildcard bins pmp20cfg = {240'b??????????????????????????????????????????1?????_??????????????????????????????????????????1?????_????????????????????????????????????????????????????????????????????????????????????01??????????_000000000000000000000000000000000000000000100000};
			wildcard bins pmp21cfg = {240'b?????????????????????????????????????????1??????_?????????????????????????????????????????1??????_??????????????????????????????????????????????????????????????????????????????????01????????????_000000000000000000000000000000000000000001000000};
			wildcard bins pmp22cfg = {240'b????????????????????????????????????????1???????_????????????????????????????????????????1???????_????????????????????????????????????????????????????????????????????????????????01??????????????_000000000000000000000000000000000000000010000000};
			wildcard bins pmp23cfg = {240'b???????????????????????????????????????1????????_???????????????????????????????????????1????????_??????????????????????????????????????????????????????????????????????????????01????????????????_000000000000000000000000000000000000000100000000};
			wildcard bins pmp24cfg = {240'b??????????????????????????????????????1?????????_??????????????????????????????????????1?????????_????????????????????????????????????????????????????????????????????????????01??????????????????_000000000000000000000000000000000000001000000000};
			wildcard bins pmp25cfg = {240'b?????????????????????????????????????1??????????_?????????????????????????????????????1??????????_??????????????????????????????????????????????????????????????????????????01????????????????????_000000000000000000000000000000000000010000000000};
			wildcard bins pmp26cfg = {240'b????????????????????????????????????1???????????_????????????????????????????????????1???????????_????????????????????????????????????????????????????????????????????????01??????????????????????_000000000000000000000000000000000000100000000000};
			wildcard bins pmp27cfg = {240'b???????????????????????????????????1????????????_???????????????????????????????????1????????????_??????????????????????????????????????????????????????????????????????01????????????????????????_000000000000000000000000000000000001000000000000};
			wildcard bins pmp28cfg = {240'b??????????????????????????????????1?????????????_??????????????????????????????????1?????????????_????????????????????????????????????????????????????????????????????01??????????????????????????_000000000000000000000000000000000010000000000000};
			wildcard bins pmp29cfg = {240'b?????????????????????????????????1??????????????_?????????????????????????????????1??????????????_??????????????????????????????????????????????????????????????????01????????????????????????????_000000000000000000000000000000000100000000000000};
			wildcard bins pmp30cfg = {240'b????????????????????????????????1???????????????_????????????????????????????????1???????????????_????????????????????????????????????????????????????????????????01??????????????????????????????_000000000000000000000000000000001000000000000000};
			wildcard bins pmp31cfg = {240'b???????????????????????????????1????????????????_???????????????????????????????1????????????????_??????????????????????????????????????????????????????????????01????????????????????????????????_000000000000000000000000000000010000000000000000};
			wildcard bins pmp32cfg = {240'b??????????????????????????????1?????????????????_??????????????????????????????1?????????????????_????????????????????????????????????????????????????????????01??????????????????????????????????_000000000000000000000000000000100000000000000000};
			wildcard bins pmp33cfg = {240'b?????????????????????????????1??????????????????_?????????????????????????????1??????????????????_??????????????????????????????????????????????????????????01????????????????????????????????????_000000000000000000000000000001000000000000000000};
			wildcard bins pmp34cfg = {240'b????????????????????????????1???????????????????_????????????????????????????1???????????????????_????????????????????????????????????????????????????????01??????????????????????????????????????_000000000000000000000000000010000000000000000000};
			wildcard bins pmp35cfg = {240'b???????????????????????????1????????????????????_???????????????????????????1????????????????????_??????????????????????????????????????????????????????01????????????????????????????????????????_000000000000000000000000000100000000000000000000};
			wildcard bins pmp36cfg = {240'b??????????????????????????1?????????????????????_??????????????????????????1?????????????????????_????????????????????????????????????????????????????01??????????????????????????????????????????_000000000000000000000000001000000000000000000000};
			wildcard bins pmp37cfg = {240'b?????????????????????????1??????????????????????_?????????????????????????1??????????????????????_??????????????????????????????????????????????????01????????????????????????????????????????????_000000000000000000000000010000000000000000000000};
			wildcard bins pmp38cfg = {240'b????????????????????????1???????????????????????_????????????????????????1???????????????????????_????????????????????????????????????????????????01??????????????????????????????????????????????_000000000000000000000000100000000000000000000000};
			wildcard bins pmp39cfg = {240'b???????????????????????1????????????????????????_???????????????????????1????????????????????????_??????????????????????????????????????????????01????????????????????????????????????????????????_000000000000000000000001000000000000000000000000};
			wildcard bins pmp40cfg = {240'b??????????????????????1?????????????????????????_??????????????????????1?????????????????????????_????????????????????????????????????????????01??????????????????????????????????????????????????_000000000000000000000010000000000000000000000000};
			wildcard bins pmp41cfg = {240'b?????????????????????1??????????????????????????_?????????????????????1??????????????????????????_??????????????????????????????????????????01????????????????????????????????????????????????????_000000000000000000000100000000000000000000000000};
			wildcard bins pmp42cfg = {240'b????????????????????1???????????????????????????_????????????????????1???????????????????????????_????????????????????????????????????????01??????????????????????????????????????????????????????_000000000000000000001000000000000000000000000000};
			wildcard bins pmp43cfg = {240'b???????????????????1????????????????????????????_???????????????????1????????????????????????????_??????????????????????????????????????01????????????????????????????????????????????????????????_000000000000000000010000000000000000000000000000};
			wildcard bins pmp44cfg = {240'b??????????????????1?????????????????????????????_??????????????????1?????????????????????????????_????????????????????????????????????01??????????????????????????????????????????????????????????_000000000000000000100000000000000000000000000000};
			wildcard bins pmp45cfg = {240'b?????????????????1??????????????????????????????_?????????????????1??????????????????????????????_??????????????????????????????????01????????????????????????????????????????????????????????????_000000000000000001000000000000000000000000000000};
			wildcard bins pmp46cfg = {240'b????????????????1???????????????????????????????_????????????????1???????????????????????????????_????????????????????????????????01??????????????????????????????????????????????????????????????_000000000000000010000000000000000000000000000000};
			wildcard bins pmp47cfg = {240'b???????????????1????????????????????????????????_???????????????1????????????????????????????????_??????????????????????????????01????????????????????????????????????????????????????????????????_000000000000000100000000000000000000000000000000};
			wildcard bins pmp48cfg = {240'b??????????????1?????????????????????????????????_??????????????1?????????????????????????????????_????????????????????????????01??????????????????????????????????????????????????????????????????_000000000000001000000000000000000000000000000000};
			wildcard bins pmp49cfg = {240'b?????????????1??????????????????????????????????_?????????????1??????????????????????????????????_??????????????????????????01????????????????????????????????????????????????????????????????????_000000000000010000000000000000000000000000000000};
			wildcard bins pmp50cfg = {240'b????????????1???????????????????????????????????_????????????1???????????????????????????????????_????????????????????????01??????????????????????????????????????????????????????????????????????_000000000000100000000000000000000000000000000000};
			wildcard bins pmp51cfg = {240'b???????????1????????????????????????????????????_???????????1????????????????????????????????????_??????????????????????01????????????????????????????????????????????????????????????????????????_000000000001000000000000000000000000000000000000};
			wildcard bins pmp52cfg = {240'b??????????1?????????????????????????????????????_??????????1?????????????????????????????????????_????????????????????01??????????????????????????????????????????????????????????????????????????_000000000010000000000000000000000000000000000000};
			wildcard bins pmp53cfg = {240'b?????????1??????????????????????????????????????_?????????1??????????????????????????????????????_??????????????????01????????????????????????????????????????????????????????????????????????????_000000000100000000000000000000000000000000000000};
			wildcard bins pmp54cfg = {240'b????????1???????????????????????????????????????_????????1???????????????????????????????????????_????????????????01??????????????????????????????????????????????????????????????????????????????_000000001000000000000000000000000000000000000000};
			wildcard bins pmp55cfg = {240'b???????1????????????????????????????????????????_???????1????????????????????????????????????????_??????????????01????????????????????????????????????????????????????????????????????????????????_000000010000000000000000000000000000000000000000};
			wildcard bins pmp56cfg = {240'b??????1?????????????????????????????????????????_??????1?????????????????????????????????????????_????????????01??????????????????????????????????????????????????????????????????????????????????_000000100000000000000000000000000000000000000000};
			wildcard bins pmp57cfg = {240'b?????1??????????????????????????????????????????_?????1??????????????????????????????????????????_??????????01????????????????????????????????????????????????????????????????????????????????????_000001000000000000000000000000000000000000000000};
			wildcard bins pmp58cfg = {240'b????1???????????????????????????????????????????_????1???????????????????????????????????????????_????????01??????????????????????????????????????????????????????????????????????????????????????_000010000000000000000000000000000000000000000000};
			wildcard bins pmp59cfg = {240'b???1????????????????????????????????????????????_???1????????????????????????????????????????????_??????01????????????????????????????????????????????????????????????????????????????????????????_000100000000000000000000000000000000000000000000};
			wildcard bins pmp61cfg = {240'b??1?????????????????????????????????????????????_??1?????????????????????????????????????????????_????01??????????????????????????????????????????????????????????????????????????????????????????_001000000000000000000000000000000000000000000000};
			wildcard bins pmp62cfg = {240'b?1??????????????????????????????????????????????_?1??????????????????????????????????????????????_??01????????????????????????????????????????????????????????????????????????????????????????????_010000000000000000000000000000000000000000000000};
			wildcard bins pmp63cfg = {240'b1???????????????????????????????????????????????_1???????????????????????????????????????????????_01??????????????????????????????????????????????????????????????????????????????????????????????_100000000000000000000000000000000000000000000000};
		}
	`endif

	rs1_val_for_pmpcfg_A: coverpoint ins.current.rs1_val {
		bins OFF = {0};
		`ifdef XLEN32
			bins TOR   = {32'b00001000000010000000100000001000};
			bins NA4   = {32'b00010000000100000001000000010000};
			bins NAPOT = {32'b00011000000110000001100000011000};
		`endif
		`ifdef XLEN64
			bins TOR   = {64'b0000100000001000000010000000100000001000000010000000100000001000};
			bins NA4   = {64'b0001000000010000000100000001000000010000000100000001000000010000};
			bins NAPOT = {64'b0001100000011000000110000001100000011000000110000001100000011000};
		`endif
	}

//-------------------------------------------------------

	// Setting the even pmpcfg to 0 and odd pmpcfg to TOR & and rotating through the 6 legal XWR values for each pair.
	pmp_entries_setup: coverpoint {pmpcfg_a[27:0], pmpcfg_l[13:0], pmpcfg_x[13:0], pmpcfg_wr[27:0]} {
		bins tor_legal_xwr = {84'b0100010001000100010001000100_10101010101010_00100010001000_0000110001000000110001000000};
	}

	overlapping_regions: coverpoint (
									 pmpaddr[13] == ((`REGIONSTART + 7*`g) >> 2) &&
									 pmpaddr[12] == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[11] == ((`REGIONSTART + 6*`g) >> 2) &&
									 pmpaddr[10] == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[9]  == ((`REGIONSTART + 5*`g) >> 2) &&
									 pmpaddr[8]  == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[7]  == ((`REGIONSTART + 4*`g) >> 2) &&
									 pmpaddr[6]  == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[5]  == ((`REGIONSTART + 3*`g) >> 2) &&
									 pmpaddr[4]  == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[3]  == ((`REGIONSTART + 2*`g) >> 2) &&
									 pmpaddr[2]  == (`REGIONSTART  >> 2)		 &&
									 pmpaddr[1]  == ((`REGIONSTART + 1*`g) >> 2) &&
									 pmpaddr[0]  == (`REGIONSTART  >> 2)
									 ) {
		bins tor_regions = {1};	// Set 1 when overlapping tor regions set up.
	}

	// Address at the end of the overlapping regions
	addr_offset_for_priority_check: coverpoint (ins.current.rs1_val+ins.current.imm) {
		bins at_end_of_region13 = {`REGIONSTART + 7*`g - 4};
		bins at_end_of_region11 = {`REGIONSTART + 6*`g - 4};
		bins at_end_of_region9  = {`REGIONSTART + 5*`g - 4};
		bins at_end_of_region7  = {`REGIONSTART + 4*`g - 4};
		bins at_end_of_region5  = {`REGIONSTART + 3*`g - 4};
		bins at_end_of_region3  = {`REGIONSTART + 2*`g - 4};
		bins at_end_of_region1  = {`REGIONSTART + 1*`g - 4};
	}

//-------------------------------------------------------

	// {TOR, OFF, TOR, OFF} and {1111, 1000, 1101, 1000}
	cfg_first_four_entries: coverpoint {pmpcfg[3],pmpcfg[2],pmpcfg[1],pmpcfg[0]} {
		bins cfg_regions = {32'h8F808D80};
	}

	first_four_pmp_entries: coverpoint (pmpaddr[0]==((`REGIONSTART)	   >> 2) &&
										pmpaddr[1]==((`REGIONSTART+`g) >> 2) &&
										pmpaddr[2]==((`REGIONSTART)	   >> 2) &&
										pmpaddr[3]==((`REGIONSTART+`g) >> 2)
										) {
		bins pmp_entries = {1};
	}

//-------------------------------------------------------

	all_pmp_entries_off: coverpoint {pmpcfg_a,pmpcfg_A[1:0]} { // Including Background Top PMP Entry
		bins PMP_OFF = {0};
	}

	// pack_pmpaddr has all the pmpaddr csrs, so when it's zero implies all pmpaddr = 0
	all_pmpaddr_zero: coverpoint pack_pmpaddr { // Including Background Top PMP Entry
		bins pmpaddr_zeros = {0};
	}

//-------------------------------------------------------

	cp_cfg_X: cross priv_mode_m, legal_lxwr, exec_instr, addr_in_region ;
	cp_cfg_R: cross priv_mode_m, legal_lxwr, read_instr, addr_in_region ;
	cp_cfg_W: cross priv_mode_m, legal_lxwr, write_instr, addr_in_region ;

	cp_cfg_X1_all: cross priv_mode_m, exec_instr, X1, addr_in_region ;
	cp_cfg_X0_all: cross priv_mode_m, exec_instr, X0, addr_in_region ;

	cp_cfg_Rw00_all: cross priv_mode_m, read_instr, RW00, addr_in_region ;
	cp_cfg_Rw10_all: cross priv_mode_m, read_instr, RW10, addr_in_region ;
	cp_cfg_Rw11_all: cross priv_mode_m, read_instr, RW11, addr_in_region ;
	cp_cfg_rW00_all: cross priv_mode_m, write_instr, RW00, addr_in_region ;
	cp_cfg_rW10_all: cross priv_mode_m, write_instr, RW10, addr_in_region ;
	cp_cfg_rW11_all: cross priv_mode_m, write_instr, RW11, addr_in_region ;

	cp_cfg_L_access_exec: cross priv_mode_m, exec_instr, RWX000, addr_in_region ;
	cp_cfg_L_access_read: cross priv_mode_m, read_instr_lw, RWX000, addr_in_region ;
	cp_cfg_L_access_write: cross priv_mode_m, write_instr_sw, RWX000, addr_in_region ;

	cp_cfg_L_modify: cross priv_mode_m, lock_checking, pmp_region, pmp_csr_to_write ;

	cp_cfg_A_all_even: cross priv_mode_m, rs1_val_for_pmpcfg_A, csrrw, legal_pmpcfg_entries_even ;
	`ifdef XLEN32
		cp_cfg_A_all_odd: cross priv_mode_m, rs1_val_for_pmpcfg_A, csrrw, legal_pmpcfg_entries_odd ;
	`endif

	cp_cfg_A_OFF_all_read : cross priv_mode_m, pmpcfgA_OFF, read_instr_lw, addr_in_region;
	cp_cfg_A_OFF_all_write : cross priv_mode_m, pmpcfgA_OFF, write_instr_sw, addr_in_region;
	cp_cfg_A_OFF_all_exec : cross priv_mode_m, pmpcfgA_OFF, exec_instr, addr_in_region;

	cp_cfg_A_napot_all: cross priv_mode_m, pmpcfgA_NAPOT, read_instr_lw, addr_offset_cp_cfg_A_napot_all;

	cp_cfg_A_napot_x : cross priv_mode_m, legal_RWX_L_NAPOT, address_offsets, exec_instr;
	cp_cfg_A_napot_r : cross priv_mode_m, legal_RWX_L_NAPOT, address_offsets, read_instr_lw;
	cp_cfg_A_napot_w : cross priv_mode_m, legal_RWX_L_NAPOT, address_offsets, write_instr_sw;

	`ifdef G_IS_0
		cp_cfg_A_NA4_all: cross priv_mode_m, pmpcfgA_NA4, read_instr_lw, addr_offset_cp_cfg_A_na4 ;

		cp_cfg_A_na4_x : cross priv_mode_m, legal_RWX_L_NA4, addr_offset_cp_cfg_A_na4, exec_instr ;
		cp_cfg_A_na4_r : cross priv_mode_m, legal_RWX_L_NA4, addr_offset_cp_cfg_A_na4, read_instr_lw ;
		cp_cfg_A_na4_w : cross priv_mode_m, legal_RWX_L_NA4, addr_offset_cp_cfg_A_na4, write_instr_sw ;
	`endif

	cp_cfg_A_tor_x : cross priv_mode_m, legal_RWX_L_TOR, address_offsets, exec_instr;
	cp_cfg_A_tor_r : cross priv_mode_m, legal_RWX_L_TOR, address_offsets, read_instr_lw;
	cp_cfg_A_tor_w : cross priv_mode_m, legal_RWX_L_TOR, address_offsets, write_instr_sw;

	cp_cfg_A_tor0_r: cross priv_mode_m, addr_offset_cp_cfg_A_tor0, pmp_addr_for_tor0,pmpcfg_for_tor0, read_instr_lw ;
	cp_cfg_A_tor0_w: cross priv_mode_m, addr_offset_cp_cfg_A_tor0, pmp_addr_for_tor0,pmpcfg_for_tor0, write_instr_sw ;
	cp_cfg_A_tor0_x: cross priv_mode_m, addr_offset_cp_cfg_A_tor0, pmp_addr_for_tor0,pmpcfg_for_tor0, exec_instr;

	cp_cfg_A_tor_all0: cross priv_mode_m, addr_for_tor_all_region0, pmpaddr_for_tor_region0, RWXL_i111_pmp0cfg, read_instr_lw;
	cp_cfg_A_tor_all1: cross priv_mode_m, addr_for_tor_all_region1, pmpaddr_for_tor_region1, RWXL_i001_pmp1cfg, read_instr_lw;
	cp_cfg_A_tor_all2: cross priv_mode_m, addr_for_tor_all_region2, pmpaddr_for_tor_region2, RWXL_i001_pmp2cfg, read_instr_lw;
	cp_cfg_A_tor_all3: cross priv_mode_m, addr_for_tor_all_region3, pmpaddr_for_tor_region3, RWXL_i001_pmp3cfg, read_instr_lw;
	cp_cfg_A_tor_all4: cross priv_mode_m, addr_for_tor_all_region4, pmpaddr_for_tor_region4, RWXL_i001_pmp4cfg, read_instr_lw;
	cp_cfg_A_tor_all5: cross priv_mode_m, addr_for_tor_all_region5, pmpaddr_for_tor_region5, RWXL_i001_pmp5cfg, read_instr_lw;
	cp_cfg_A_tor_all6: cross priv_mode_m, addr_for_tor_all_region6, pmpaddr_for_tor_region6, RWXL_i001_pmp6cfg, read_instr_lw;
	cp_cfg_A_tor_all7: cross priv_mode_m, addr_for_tor_all_region7, pmpaddr_for_tor_region7, RWXL_i001_pmp7cfg, read_instr_lw;
	cp_cfg_A_tor_all8: cross priv_mode_m, addr_for_tor_all_region8, pmpaddr_for_tor_region8, RWXL_i001_pmp8cfg, read_instr_lw;
	cp_cfg_A_tor_all9: cross priv_mode_m, addr_for_tor_all_region9, pmpaddr_for_tor_region9, RWXL_i001_pmp9cfg, read_instr_lw;
	cp_cfg_A_tor_all10: cross priv_mode_m, addr_for_tor_all_region10, pmpaddr_for_tor_region10, RWXL_i001_pmp10cfg, read_instr_lw;
	cp_cfg_A_tor_all11: cross priv_mode_m, addr_for_tor_all_region11, pmpaddr_for_tor_region11, RWXL_i001_pmp11cfg, read_instr_lw;
	cp_cfg_A_tor_all12: cross priv_mode_m, addr_for_tor_all_region12, pmpaddr_for_tor_region12, RWXL_i001_pmp12cfg, read_instr_lw;
	cp_cfg_A_tor_all13: cross priv_mode_m, addr_for_tor_all_region13, pmpaddr_for_tor_region13, RWXL_i001_pmp13cfg, read_instr_lw;
	cp_cfg_A_tor_all14: cross priv_mode_m, addr_for_tor_all_region14, pmpaddr_for_tor_region14, RWXL_i001_pmp14cfg, read_instr_lw;

	cp_cfg_A_tor_bot_L0_x: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L0, pmp_addr_for_tor_bot, exec_instr;
	cp_cfg_A_tor_bot_L0_w: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L0, pmp_addr_for_tor_bot, write_instr_sw;
	cp_cfg_A_tor_bot_L0_r: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L0, pmp_addr_for_tor_bot, read_instr_lw;

	cp_cfg_A_tor_bot_L1_x: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L1, pmp_addr_for_tor_bot, exec_instr;
	cp_cfg_A_tor_bot_L1_w: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L1, pmp_addr_for_tor_bot, write_instr_sw;
	cp_cfg_A_tor_bot_L1_r: cross priv_mode_m, addr_for_tor_bot, pmpcfg_tor_bot_L1, pmp_addr_for_tor_bot, read_instr_lw;

	cp_cfg_A_tor_nonoverlap1_x: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap1, exec_instr;
	cp_cfg_A_tor_nonoverlap1_w: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap1, write_instr_sw;
	cp_cfg_A_tor_nonoverlap1_r: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap1, read_instr_lw;

	cp_cfg_A_tor_nonoverlap2_x: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap2, exec_instr;
	cp_cfg_A_tor_nonoverlap2_w: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap2, write_instr_sw;
	cp_cfg_A_tor_nonoverlap2_r: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap2, read_instr_lw;

	cp_cfg_A_tor_nonoverlap3_x: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap3, exec_instr;
	cp_cfg_A_tor_nonoverlap3_w: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap3, write_instr_sw;
	cp_cfg_A_tor_nonoverlap3_r: cross priv_mode_m, addr_for_tor_nonoverlap, pmpcfg_tor_nonoverlap, pmp_addr_for_tor_nonoverlap3, read_instr_lw;

	cp_pmpaddr_walk: cross priv_mode_m, cp_walk_rs1, csrrw, legal_pmpaddr_entries ;
	cp_pmpcfg_walk: cross priv_mode_m, cp_walk_rs1, csrrw, legal_pmpcfg_entries_even ;
	`ifdef XLEN32
		// Will throw illegal instruction when XLEN = 64.
		cp_pmpcfg_zero: cross priv_mode_m, cp_zero_rs1, csrrw, legal_pmpcfg_entries_odd ;
	`endif

	`ifdef PMP_64
		cp_pmp64_write: cross priv_mode_m, write_instr_sw, pmp64;
		cp_pmp64_read: cross priv_mode_m, read_instr_lw, pmp64;
	`endif

	cp_priority_lw: cross priv_mode_m, pmp_entries_setup, overlapping_regions, addr_offset_for_priority_check, read_instr_lw ;
	cp_priority_sw: cross priv_mode_m, pmp_entries_setup, overlapping_regions, addr_offset_for_priority_check, write_instr_sw ;
	cp_priority_jalr: cross priv_mode_m, pmp_entries_setup, overlapping_regions, addr_offset_for_priority_check, exec_instr ;

	cp_priority_off_lw: cross priv_mode_m, cfg_first_four_entries, first_four_pmp_entries, read_instr_lw ;
	cp_priority_off_sw: cross priv_mode_m, cfg_first_four_entries, first_four_pmp_entries, write_instr_sw ;
	cp_priority_off_jalr: cross priv_mode_m, cfg_first_four_entries, first_four_pmp_entries, exec_instr ;

	cp_none_lw: cross priv_mode_m, all_pmp_entries_off, all_pmpaddr_zero, read_instr_lw ;
	cp_none_sw: cross priv_mode_m, all_pmp_entries_off, all_pmpaddr_zero, write_instr_sw ;
	cp_none_jalr: cross priv_mode_m, all_pmp_entries_off, all_pmpaddr_zero, exec_instr ;

	// For cp_grain, writing and reading from pmpaddr0 and pmpcfg0 is a part of the test, even though it is
	// too dificult to check with the coverpoint. Below is the snippet of the code

	/*li t0, 8'b00011111
	li t1, 8'b00000111
	csrw pmpcfg0, t0 #pmpcfg0.A = NAPOT
	li t0, {0/1s/checkerboard}
	csrw pmpaddr0, t0 # pmpaddr0 = value under test
	csrr t2, pmpaddr0
	SIGUPD(t2) # read back pmpaddr0, which should have G-1 trailing 1s
	csrw pmpcfg0, t1 # pmpcfg0.A = OFF
	csrr t2, pmpaddr0
	SIGUPD(t2) # read back pmpaddr0, which should have G trailing 0s*/
	`ifndef G_IS_0
		cp_grain_OFF_to_OFF : cross priv_mode_m, pmpcfg0_A_mode_was_OFF, pmpcfg0_A_mode_is_OFF ;
		cp_grain_OFF_to_NAPOT : cross priv_mode_m, pmpcfg0_A_mode_was_OFF, pmpcfg0_A_mode_is_NAPOT ;
		cp_grain_OFF_to_TOR : cross priv_mode_m, pmpcfg0_A_mode_was_OFF, pmpcfg0_A_mode_is_TOR ;
		cp_grain_NAPOT_to_OFF : cross priv_mode_m, pmpcfg0_A_mode_was_NAPOT, pmpcfg0_A_mode_is_OFF ;
		cp_grain_NAPOT_to_NAPOT : cross priv_mode_m, pmpcfg0_A_mode_was_NAPOT, pmpcfg0_A_mode_is_NAPOT ;
		cp_grain_NAPOT_to_TOR : cross priv_mode_m, pmpcfg0_A_mode_was_NAPOT, pmpcfg0_A_mode_is_TOR ;
	`endif

	cp_grain_check: cross priv_mode_m, pmpcfg_for_cp_grain_check, pmpaddr0_for_cp_grain_check, csrrw_to_pmpaddr0, csrr_to_pmpaddr0;

	//crosses boundary for napot region at the start of the region.
	cp_misaligned_napot_start_r: cross priv_mode_m, pmpaddr_for_napot_misaligned, pmpcfg_for_napot_misaligned, addr_for_misaligned_straddling_start, read_instr_for_misaligned;
	cp_misaligned_napot_start_w: cross priv_mode_m, pmpaddr_for_napot_misaligned, pmpcfg_for_napot_misaligned, addr_for_misaligned_straddling_start, write_instr_for_misaligned;

	//crosses boundary for napot region at the end of the region.
	cp_misaligned_napot_end_r: cross priv_mode_m, pmpaddr_for_napot_misaligned, pmpcfg_for_napot_misaligned, addr_for_misaligned_straddling_end, read_instr_for_misaligned;
	cp_misaligned_napot_end_w: cross priv_mode_m, pmpaddr_for_napot_misaligned, pmpcfg_for_napot_misaligned, addr_for_misaligned_straddling_end, write_instr_for_misaligned;

	cp_misaligned_tor_start_r: cross priv_mode_m, pmpaddr_for_tor_misaligned, pmpcfg_for_tor_misaligned, addr_for_misaligned_straddling_start, read_instr_for_misaligned;
	cp_misaligned_tor_start_w: cross priv_mode_m, pmpaddr_for_tor_misaligned, pmpcfg_for_tor_misaligned, addr_for_misaligned_straddling_start, write_instr_for_misaligned;

	cp_misaligned_tor_end_r: cross priv_mode_m, pmpaddr_for_tor_misaligned, pmpcfg_for_tor_misaligned, addr_for_misaligned_straddling_end, read_instr_for_misaligned;
	cp_misaligned_tor_end_w: cross priv_mode_m, pmpaddr_for_tor_misaligned, pmpcfg_for_tor_misaligned, addr_for_misaligned_straddling_end, write_instr_for_misaligned;

	cp_misaligned_off_start_r: cross priv_mode_m, pmpaddr_for_off_misaligned, pmpcfg_for_off_misaligned, addr_for_misaligned_straddling_start, read_instr_for_misaligned;
	cp_misaligned_off_start_w: cross priv_mode_m, pmpaddr_for_off_misaligned, pmpcfg_for_off_misaligned, addr_for_misaligned_straddling_start, write_instr_for_misaligned;

	cp_misaligned_off_end_r: cross priv_mode_m, pmpaddr_for_off_misaligned, pmpcfg_for_off_misaligned, addr_for_misaligned_straddling_end, read_instr_for_misaligned;
	cp_misaligned_off_end_w: cross priv_mode_m, pmpaddr_for_off_misaligned, pmpcfg_for_off_misaligned, addr_for_misaligned_straddling_end, write_instr_for_misaligned;

	`ifdef G_IS_0
		cp_misaligned_na4_start_r: cross priv_mode_m, pmpaddr_for_na4_misaligned, pmpcfg_for_na4_misaligned, addr_for_na4_misaligned_straddling_start, read_instr_for_misaligned;
		cp_misaligned_na4_start_w: cross priv_mode_m, pmpaddr_for_na4_misaligned, pmpcfg_for_na4_misaligned, addr_for_na4_misaligned_straddling_start, write_instr_for_misaligned;

		cp_misaligned_na4_end_r: cross priv_mode_m, pmpaddr_for_na4_misaligned, pmpcfg_for_na4_misaligned, addr_for_na4_misaligned_straddling_end, read_instr_for_misaligned;
		cp_misaligned_na4_end_w: cross priv_mode_m, pmpaddr_for_na4_misaligned, pmpcfg_for_na4_misaligned, addr_for_na4_misaligned_straddling_end, write_instr_for_misaligned;
	`endif

  `ifdef XLEN64
		`ifdef G_IS_0
			pmpaddr_for_na4_even: coverpoint {pmpaddr[0]} {
				bins address_even = {`NON_STANDARD_REGION};
			}

			pmpaddr_for_na4_odd: coverpoint {pmpaddr[1]} {
				bins address_odd = {`NON_STANDARD_REGION+4};
			}

			pmpcfg_na4_lxwr_even: coverpoint pmpcfg[0] {
				bins locked_na4_region = {8'b10010111};
			}

			pmpcfg_na4_lxwr_odd: coverpoint pmpcfg[1] {
				bins locked_na4_region = {8'b10010111};
			}

			addr_for_na4: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {`NON_STANDARD_REGION<<2};
			}

			pmpaddr_for_tor_even: coverpoint {pmpaddr[1],pmpaddr[0]}  {
				bins four_byte_tor = {`NON_STANDARD_REGION+1,`NON_STANDARD_REGION};
			}

			pmpaddr_for_tor_odd: coverpoint {pmpaddr[3],pmpaddr[2]}  {
				bins four_byte_tor = {`NON_STANDARD_REGION+4,`NON_STANDARD_REGION+3};
			}

			addr_for_tor_odd: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {(`NON_STANDARD_REGION<<2)+8};
			}

			addr_for_tor_even: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {`NON_STANDARD_REGION<<2};
			}

			pmpcfg_tor_lxwr_even: coverpoint {pmpcfg[1],pmpcfg[0]} {
				bins locked_tor_region = {16'b10001111_00000111};
			}

			pmpcfg_tor_lxwr_odd: coverpoint {pmpcfg[3],pmpcfg[2]} {
				bins locked_tor_region = {16'b10001111_00000111};
			}

			pmpaddr_for_double_tor: coverpoint {pmpaddr[5],pmpaddr[4],pmpaddr[3]}  {
				bins byte_double_tor = {`NON_STANDARD_REGION+6,`NON_STANDARD_REGION+5,`NON_STANDARD_REGION+4};
			}

			pmpcfg_double_tor_lxwr: coverpoint {pmpcfg[5],pmpcfg[4]}  {
				bins locked_tor_region = {16'b1000111110001111};
			}

			addr_for_tor_double: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {(`NON_STANDARD_REGION<<2)+16};
			}

			pmpcfg_for_na4_wrap: coverpoint pmpcfg[0] {
				bins na4_wrap_locked = {8'b10010111};
				bins na4_wrap_unlocked = {8'b00010111};
			}

			addr_for_na4_wrap: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {(`NON_STANDARD_REGION<<2)-2};
			}

			pmpaddr_for_tor_wrap: coverpoint {pmpaddr[1],pmpaddr[0]}  {
				bins four_byte_tor = {`NON_STANDARD_REGION+1,`NON_STANDARD_REGION};
			}

			pmpcfg_for_tor_wrap: coverpoint {pmpcfg[1],pmpcfg[0]} {
				bins tor_wrap_locked = {16'b10001111_10001111};
				bins tor_wrap_unlocked = {16'b00001111_00001111};
			}

			addr_for_tor_wrap: coverpoint (ins.current.rs1_val + ins.current.imm) {
				bins address_to_access = {(`NON_STANDARD_REGION<<2)-2};
			}

			read_instr_ld: coverpoint ins.current.insn {
    			wildcard bins ld = {32'b?????????????????_011?????_0000011};
			}

			write_instr_sd: coverpoint ins.current.insn {
				wildcard bins sd = {32'b?????????????????_011?????_0100011};
			}

			cp_na4_boundary_ld_even: cross priv_mode_m, pmpaddr_for_na4_even, pmpcfg_na4_lxwr_even, read_instr_ld, addr_for_na4 ;
			cp_na4_boundary_ld_odd: cross priv_mode_m, pmpaddr_for_na4_odd, pmpcfg_na4_lxwr_odd, read_instr_ld, addr_for_na4 ;

			cp_na4_boundary_sd_even: cross priv_mode_m, pmpaddr_for_na4_even, pmpcfg_na4_lxwr_even, write_instr_sd, addr_for_na4  ;
			cp_na4_boundary_sd_odd: cross priv_mode_m, pmpaddr_for_na4_odd, pmpcfg_na4_lxwr_odd, write_instr_sd, addr_for_na4  ;

			cp_tor_boundary_ld_even: cross priv_mode_m, pmpaddr_for_tor_even, pmpcfg_tor_lxwr_even, read_instr_ld, addr_for_tor_even ;
			cp_tor_boundary_ld_odd: cross priv_mode_m, pmpaddr_for_tor_odd, pmpcfg_tor_lxwr_odd, read_instr_ld, addr_for_tor_odd ;

			cp_tor_boundary_sd_even: cross priv_mode_m, pmpaddr_for_tor_even, pmpcfg_tor_lxwr_even, write_instr_sd, addr_for_tor_even  ;
			cp_tor_boundary_sd_odd: cross priv_mode_m, pmpaddr_for_tor_odd, pmpcfg_tor_lxwr_odd, write_instr_sd, addr_for_tor_odd  ;

			cp_tor_doubleregionfail_ld: cross priv_mode_m, pmpaddr_for_double_tor, pmpcfg_double_tor_lxwr, read_instr_ld, addr_for_tor_double ;
			cp_tor_doubleregionfail_sd: cross priv_mode_m, pmpaddr_for_double_tor, pmpcfg_double_tor_lxwr, write_instr_sd, addr_for_tor_double  ;

			cp_misaligned_na4_wrap_ld: cross priv_mode_m, pmpaddr_for_na4_even, pmpcfg_for_na4_wrap, read_instr_ld, addr_for_na4_wrap ;
			cp_misaligned_na4_wrap_sd: cross priv_mode_m, pmpaddr_for_na4_even, pmpcfg_for_na4_wrap, write_instr_sd, addr_for_na4_wrap ;

			cp_misaligned_tor_wrap_ld: cross priv_mode_m, pmpaddr_for_tor_wrap, pmpcfg_for_tor_wrap, read_instr_ld, addr_for_tor_wrap ;
			cp_misaligned_tor_wrap_sd: cross priv_mode_m, pmpaddr_for_tor_wrap, pmpcfg_for_tor_wrap, write_instr_sd, addr_for_tor_wrap ;
		`endif
	`endif

endgroup

function void pmpm_sample(int hart, int issue, ins_t ins);

	logic [7:0] pmpcfg [63:0];
	logic [XLEN-1:0] pmpaddr [62:0];
	logic [16*XLEN-1:0] pack_pmpaddr;
	logic [29:0] pmpcfg_wr, pmpcfg_a;			// for first 15 Regions
	logic [95:0] pmpcfg_WR, pmpcfg_A;			// for next 48 Regions
	logic [14:0] pmpcfg_x, pmpcfg_l, pmp_hit;   // for first 15 Regions
	logic [47:0] pmpcfg_X, pmpcfg_L, pmp_HIT;   // for next 48 Regions

	`ifdef XLEN32
	    // Each pmpcfg CSR holds 4 region configs in 32-bit (4x 8-bit)
    	for (int i = 0; i < 16; i++) begin
    	    logic [31:0] cfg_word = ins.current.csr[12'h3A0 + i];
    	    pmpcfg[i*4 + 0] = cfg_word[7:0];
    	    pmpcfg[i*4 + 1] = cfg_word[15:8];
    	    pmpcfg[i*4 + 2] = cfg_word[23:16];
    	    pmpcfg[i*4 + 3] = cfg_word[31:24];
    	end
	`elsif XLEN64
	    // Each pmpcfg CSR holds 8 region configs in 64-bit (8x 8-bit)
		for (int i = 0; i < 8; i++) begin
		    logic [63:0] cfg_word = ins.current.csr[12'h3A0 + 2*i];
		    pmpcfg[i*8 + 0] = cfg_word[7:0];
		    pmpcfg[i*8 + 1] = cfg_word[15:8];
		    pmpcfg[i*8 + 2] = cfg_word[23:16];
		    pmpcfg[i*8 + 3] = cfg_word[31:24];
		    pmpcfg[i*8 + 4] = cfg_word[39:32];
		    pmpcfg[i*8 + 5] = cfg_word[47:40];
		    pmpcfg[i*8 + 6] = cfg_word[55:48];
		    pmpcfg[i*8 + 7] = cfg_word[63:56];
		end
	`endif

	for (int j = 0; j < 63; j++) begin
		pmpaddr[j] = ins.current.csr[12'h3B0 + j];
	end

	for (int k = 0; k < 15; k++) begin  // Check for first 15 PMP regions
		pmp_hit[k] = (pmpaddr[k] == `STANDARD_REGION) || (pmpaddr[k] == `NON_STANDARD_REGION);
	end

	for (int k = 15; k < 63; k++) begin				// for next 48 regions
		pmp_HIT[k-15] = (pmpaddr[k] == `STANDARD_REGION);
	end

	pack_pmpaddr = {  ins.current.csr[12'h3BF]
					 ,ins.current.csr[12'h3BE]
					 ,ins.current.csr[12'h3BD]
					 ,ins.current.csr[12'h3BC]
					 ,ins.current.csr[12'h3BB]
					 ,ins.current.csr[12'h3BA]
					 ,ins.current.csr[12'h3B9]
					 ,ins.current.csr[12'h3B8]
					 ,ins.current.csr[12'h3B7]
					 ,ins.current.csr[12'h3B6]
					 ,ins.current.csr[12'h3B5]
					 ,ins.current.csr[12'h3B4]
					 ,ins.current.csr[12'h3B3]
					 ,ins.current.csr[12'h3B2]
					 ,ins.current.csr[12'h3B1]
					 ,ins.current.csr[12'h3B0]
					};

	`ifdef XLEN32
		pmpcfg_wr = {
					ins.current.csr[12'h3A3][17:16],
					ins.current.csr[12'h3A3][9:8],
					ins.current.csr[12'h3A3][1:0],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A1][25:24],
					ins.current.csr[12'h3A1][17:16],
					ins.current.csr[12'h3A1][9:8],
					ins.current.csr[12'h3A1][1:0],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_wr = {
					ins.current.csr[12'h3A2][49:48],
					ins.current.csr[12'h3A2][41:40],
					ins.current.csr[12'h3A2][33:32],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A0][57:56],
					ins.current.csr[12'h3A0][49:48],
					ins.current.csr[12'h3A0][41:40],
					ins.current.csr[12'h3A0][33:32],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_WR = {
					ins.current.csr[12'h3AF][17:16],
					ins.current.csr[12'h3AF][9:8],
					ins.current.csr[12'h3AF][1:0],
					ins.current.csr[12'h3AE][25:24],
					ins.current.csr[12'h3AE][17:16],
					ins.current.csr[12'h3AE][9:8],
					ins.current.csr[12'h3AE][1:0],
					ins.current.csr[12'h3AD][25:24],
					ins.current.csr[12'h3AD][17:16],
					ins.current.csr[12'h3AD][9:8],
					ins.current.csr[12'h3AD][1:0],
					ins.current.csr[12'h3AC][25:24],
					ins.current.csr[12'h3AC][17:16],
					ins.current.csr[12'h3AC][9:8],
					ins.current.csr[12'h3AC][1:0],
					ins.current.csr[12'h3AB][25:24],
					ins.current.csr[12'h3AB][17:16],
					ins.current.csr[12'h3AB][9:8],
					ins.current.csr[12'h3AB][1:0],
					ins.current.csr[12'h3AA][25:24],
					ins.current.csr[12'h3AA][17:16],
					ins.current.csr[12'h3AA][9:8],
					ins.current.csr[12'h3AA][1:0],
					ins.current.csr[12'h3A9][25:24],
					ins.current.csr[12'h3A9][17:16],
					ins.current.csr[12'h3A9][9:8],
					ins.current.csr[12'h3A9][1:0],
					ins.current.csr[12'h3A8][25:24],
					ins.current.csr[12'h3A8][17:16],
					ins.current.csr[12'h3A8][9:8],
					ins.current.csr[12'h3A8][1:0],
					ins.current.csr[12'h3A7][25:24],
					ins.current.csr[12'h3A7][17:16],
					ins.current.csr[12'h3A7][9:8],
					ins.current.csr[12'h3A7][1:0],
					ins.current.csr[12'h3A6][25:24],
					ins.current.csr[12'h3A6][17:16],
					ins.current.csr[12'h3A6][9:8],
					ins.current.csr[12'h3A6][1:0],
					ins.current.csr[12'h3A5][25:24],
					ins.current.csr[12'h3A5][17:16],
					ins.current.csr[12'h3A5][9:8],
					ins.current.csr[12'h3A5][1:0],
					ins.current.csr[12'h3A4][25:24],
					ins.current.csr[12'h3A4][17:16],
					ins.current.csr[12'h3A4][9:8],
					ins.current.csr[12'h3A4][1:0],
					ins.current.csr[12'h3A3][25:24]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_WR = {
					ins.current.csr[12'h3AE][49:48],
					ins.current.csr[12'h3AE][41:40],
					ins.current.csr[12'h3AE][33:32],
					ins.current.csr[12'h3AE][25:24],
					ins.current.csr[12'h3AE][17:16],
					ins.current.csr[12'h3AE][9:8],
					ins.current.csr[12'h3AE][1:0],
					ins.current.csr[12'h3AC][57:56],
					ins.current.csr[12'h3AC][49:48],
					ins.current.csr[12'h3AC][41:40],
					ins.current.csr[12'h3AC][33:32],
					ins.current.csr[12'h3AC][25:24],
					ins.current.csr[12'h3AC][17:16],
					ins.current.csr[12'h3AC][9:8],
					ins.current.csr[12'h3AC][1:0],
					ins.current.csr[12'h3AA][57:56],
					ins.current.csr[12'h3AA][49:48],
					ins.current.csr[12'h3AA][41:40],
					ins.current.csr[12'h3AA][33:32],
					ins.current.csr[12'h3AA][25:24],
					ins.current.csr[12'h3AA][17:16],
					ins.current.csr[12'h3AA][9:8],
					ins.current.csr[12'h3AA][1:0],
					ins.current.csr[12'h3A8][57:56],
					ins.current.csr[12'h3A8][49:48],
					ins.current.csr[12'h3A8][41:40],
					ins.current.csr[12'h3A8][33:32],
					ins.current.csr[12'h3A8][25:24],
					ins.current.csr[12'h3A8][17:16],
					ins.current.csr[12'h3A8][9:8],
					ins.current.csr[12'h3A8][1:0],
					ins.current.csr[12'h3A6][57:56],
					ins.current.csr[12'h3A6][49:48],
					ins.current.csr[12'h3A6][41:40],
					ins.current.csr[12'h3A6][33:32],
					ins.current.csr[12'h3A6][25:24],
					ins.current.csr[12'h3A6][17:16],
					ins.current.csr[12'h3A6][9:8],
					ins.current.csr[12'h3A6][1:0],
					ins.current.csr[12'h3A4][57:56],
					ins.current.csr[12'h3A4][49:48],
					ins.current.csr[12'h3A4][41:40],
					ins.current.csr[12'h3A4][33:32],
					ins.current.csr[12'h3A4][25:24],
					ins.current.csr[12'h3A4][17:16],
					ins.current.csr[12'h3A4][9:8],
					ins.current.csr[12'h3A4][1:0],
					ins.current.csr[12'h3A2][57:56]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_X =  {
					ins.current.csr[12'h3AF][18],
					ins.current.csr[12'h3AF][10],
					ins.current.csr[12'h3AF][2],
					ins.current.csr[12'h3AE][26],
					ins.current.csr[12'h3AE][18],
					ins.current.csr[12'h3AE][10],
					ins.current.csr[12'h3AE][2],
					ins.current.csr[12'h3AD][26],
					ins.current.csr[12'h3AD][18],
					ins.current.csr[12'h3AD][10],
					ins.current.csr[12'h3AD][2],
					ins.current.csr[12'h3AC][26],
					ins.current.csr[12'h3AC][18],
					ins.current.csr[12'h3AC][10],
					ins.current.csr[12'h3AC][2],
					ins.current.csr[12'h3AB][26],
					ins.current.csr[12'h3AB][18],
					ins.current.csr[12'h3AB][10],
					ins.current.csr[12'h3AB][2],
					ins.current.csr[12'h3AA][26],
					ins.current.csr[12'h3AA][18],
					ins.current.csr[12'h3AA][10],
					ins.current.csr[12'h3AA][2],
					ins.current.csr[12'h3A9][26],
					ins.current.csr[12'h3A9][18],
					ins.current.csr[12'h3A9][10],
					ins.current.csr[12'h3A9][2],
					ins.current.csr[12'h3A8][26],
					ins.current.csr[12'h3A8][18],
					ins.current.csr[12'h3A8][10],
					ins.current.csr[12'h3A8][2],
					ins.current.csr[12'h3A7][26],
					ins.current.csr[12'h3A7][18],
					ins.current.csr[12'h3A7][10],
					ins.current.csr[12'h3A7][2],
					ins.current.csr[12'h3A6][26],
					ins.current.csr[12'h3A6][18],
					ins.current.csr[12'h3A6][10],
					ins.current.csr[12'h3A6][2],
					ins.current.csr[12'h3A5][26],
					ins.current.csr[12'h3A5][18],
					ins.current.csr[12'h3A5][10],
					ins.current.csr[12'h3A5][2],
					ins.current.csr[12'h3A4][26],
					ins.current.csr[12'h3A4][18],
					ins.current.csr[12'h3A4][10],
					ins.current.csr[12'h3A4][2],
					ins.current.csr[12'h3A3][18]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_X =  {
					ins.current.csr[12'h3AE][50],
					ins.current.csr[12'h3AE][42],
					ins.current.csr[12'h3AE][34],
					ins.current.csr[12'h3AE][26],
					ins.current.csr[12'h3AE][18],
					ins.current.csr[12'h3AE][10],
					ins.current.csr[12'h3AE][2],
					ins.current.csr[12'h3AC][58],
					ins.current.csr[12'h3AC][50],
					ins.current.csr[12'h3AC][42],
					ins.current.csr[12'h3AC][34],
					ins.current.csr[12'h3AC][26],
					ins.current.csr[12'h3AC][18],
					ins.current.csr[12'h3AC][10],
					ins.current.csr[12'h3AC][2],
					ins.current.csr[12'h3AA][58],
					ins.current.csr[12'h3AA][50],
					ins.current.csr[12'h3AA][42],
					ins.current.csr[12'h3AA][34],
					ins.current.csr[12'h3AA][26],
					ins.current.csr[12'h3AA][18],
					ins.current.csr[12'h3AA][10],
					ins.current.csr[12'h3AA][2],
					ins.current.csr[12'h3A8][58],
					ins.current.csr[12'h3A8][50],
					ins.current.csr[12'h3A8][42],
					ins.current.csr[12'h3A8][34],
					ins.current.csr[12'h3A8][26],
					ins.current.csr[12'h3A8][18],
					ins.current.csr[12'h3A8][10],
					ins.current.csr[12'h3A8][2],
					ins.current.csr[12'h3A6][58],
					ins.current.csr[12'h3A6][50],
					ins.current.csr[12'h3A6][42],
					ins.current.csr[12'h3A6][34],
					ins.current.csr[12'h3A6][26],
					ins.current.csr[12'h3A6][18],
					ins.current.csr[12'h3A6][10],
					ins.current.csr[12'h3A6][2],
					ins.current.csr[12'h3A4][58],
					ins.current.csr[12'h3A4][50],
					ins.current.csr[12'h3A4][42],
					ins.current.csr[12'h3A4][34],
					ins.current.csr[12'h3A4][26],
					ins.current.csr[12'h3A4][18],
					ins.current.csr[12'h3A4][10],
					ins.current.csr[12'h3A4][2],
					ins.current.csr[12'h3A2][58]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_x =  {
					ins.current.csr[12'h3A3][18],
					ins.current.csr[12'h3A3][10],
					ins.current.csr[12'h3A3][2],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A1][26],
					ins.current.csr[12'h3A1][18],
					ins.current.csr[12'h3A1][10],
					ins.current.csr[12'h3A1][2],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_x =  {
					ins.current.csr[12'h3A2][50],
					ins.current.csr[12'h3A2][42],
					ins.current.csr[12'h3A2][34],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A0][58],
					ins.current.csr[12'h3A0][50],
					ins.current.csr[12'h3A0][42],
					ins.current.csr[12'h3A0][34],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_a =  {
					ins.current.csr[12'h3A3][20:19],
					ins.current.csr[12'h3A3][12:11],
					ins.current.csr[12'h3A3][4:3],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A1][28:27],
					ins.current.csr[12'h3A1][20:19],
					ins.current.csr[12'h3A1][12:11],
					ins.current.csr[12'h3A1][4:3],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_a =  {
					ins.current.csr[12'h3A2][52:51],
					ins.current.csr[12'h3A2][44:43],
					ins.current.csr[12'h3A2][36:35],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A0][60:59],
					ins.current.csr[12'h3A0][52:51],
					ins.current.csr[12'h3A0][44:43],
					ins.current.csr[12'h3A0][36:35],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_A =  {
					ins.current.csr[12'h3AF][20:19],
					ins.current.csr[12'h3AF][12:11],
					ins.current.csr[12'h3AF][4:3],
					ins.current.csr[12'h3AE][28:27],
					ins.current.csr[12'h3AE][20:19],
					ins.current.csr[12'h3AE][12:11],
					ins.current.csr[12'h3AE][4:3],
					ins.current.csr[12'h3AD][28:27],
					ins.current.csr[12'h3AD][20:19],
					ins.current.csr[12'h3AD][12:11],
					ins.current.csr[12'h3AD][4:3],
					ins.current.csr[12'h3AC][28:27],
					ins.current.csr[12'h3AC][20:19],
					ins.current.csr[12'h3AC][12:11],
					ins.current.csr[12'h3AC][4:3],
					ins.current.csr[12'h3AB][28:27],
					ins.current.csr[12'h3AB][20:19],
					ins.current.csr[12'h3AB][12:11],
					ins.current.csr[12'h3AB][4:3],
					ins.current.csr[12'h3AA][28:27],
					ins.current.csr[12'h3AA][20:19],
					ins.current.csr[12'h3AA][12:11],
					ins.current.csr[12'h3AA][4:3],
					ins.current.csr[12'h3A9][28:27],
					ins.current.csr[12'h3A9][20:19],
					ins.current.csr[12'h3A9][12:11],
					ins.current.csr[12'h3A9][4:3],
					ins.current.csr[12'h3A8][28:27],
					ins.current.csr[12'h3A8][20:19],
					ins.current.csr[12'h3A8][12:11],
					ins.current.csr[12'h3A8][4:3],
					ins.current.csr[12'h3A7][28:27],
					ins.current.csr[12'h3A7][20:19],
					ins.current.csr[12'h3A7][12:11],
					ins.current.csr[12'h3A7][4:3],
					ins.current.csr[12'h3A6][28:27],
					ins.current.csr[12'h3A6][20:19],
					ins.current.csr[12'h3A6][12:11],
					ins.current.csr[12'h3A6][4:3],
					ins.current.csr[12'h3A5][28:27],
					ins.current.csr[12'h3A5][20:19],
					ins.current.csr[12'h3A5][12:11],
					ins.current.csr[12'h3A5][4:3],
					ins.current.csr[12'h3A4][28:27],
					ins.current.csr[12'h3A4][20:19],
					ins.current.csr[12'h3A4][12:11],
					ins.current.csr[12'h3A4][4:3],
					ins.current.csr[12'h3A3][28:27]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_A =  {
					ins.current.csr[12'h3AE][52:51],
					ins.current.csr[12'h3AE][44:43],
					ins.current.csr[12'h3AE][36:35],
					ins.current.csr[12'h3AE][28:27],
					ins.current.csr[12'h3AE][20:19],
					ins.current.csr[12'h3AE][12:11],
					ins.current.csr[12'h3AE][4:3],
					ins.current.csr[12'h3AC][60:59],
					ins.current.csr[12'h3AC][52:51],
					ins.current.csr[12'h3AC][44:43],
					ins.current.csr[12'h3AC][36:35],
					ins.current.csr[12'h3AC][28:27],
					ins.current.csr[12'h3AC][20:19],
					ins.current.csr[12'h3AC][12:11],
					ins.current.csr[12'h3AC][4:3],
					ins.current.csr[12'h3AA][60:59],
					ins.current.csr[12'h3AA][52:51],
					ins.current.csr[12'h3AA][44:43],
					ins.current.csr[12'h3AA][36:35],
					ins.current.csr[12'h3AA][28:27],
					ins.current.csr[12'h3AA][20:19],
					ins.current.csr[12'h3AA][12:11],
					ins.current.csr[12'h3AA][4:3],
					ins.current.csr[12'h3A8][60:59],
					ins.current.csr[12'h3A8][52:51],
					ins.current.csr[12'h3A8][44:43],
					ins.current.csr[12'h3A8][36:35],
					ins.current.csr[12'h3A8][28:27],
					ins.current.csr[12'h3A8][20:19],
					ins.current.csr[12'h3A8][12:11],
					ins.current.csr[12'h3A8][4:3],
					ins.current.csr[12'h3A6][60:59],
					ins.current.csr[12'h3A6][52:51],
					ins.current.csr[12'h3A6][44:43],
					ins.current.csr[12'h3A6][36:35],
					ins.current.csr[12'h3A6][28:27],
					ins.current.csr[12'h3A6][20:19],
					ins.current.csr[12'h3A6][12:11],
					ins.current.csr[12'h3A6][4:3],
					ins.current.csr[12'h3A4][60:59],
					ins.current.csr[12'h3A4][52:51],
					ins.current.csr[12'h3A4][44:43],
					ins.current.csr[12'h3A4][36:35],
					ins.current.csr[12'h3A4][28:27],
					ins.current.csr[12'h3A4][20:19],
					ins.current.csr[12'h3A4][12:11],
					ins.current.csr[12'h3A4][4:3],
					ins.current.csr[12'h3A2][60:59]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_L =  {
					ins.current.csr[12'h3AF][23],
					ins.current.csr[12'h3AF][15],
					ins.current.csr[12'h3AF][7],
					ins.current.csr[12'h3AD][31],
					ins.current.csr[12'h3AD][23],
					ins.current.csr[12'h3AD][15],
					ins.current.csr[12'h3AD][7],
					ins.current.csr[12'h3AD][31],
					ins.current.csr[12'h3AD][23],
					ins.current.csr[12'h3AD][15],
					ins.current.csr[12'h3AD][7],
					ins.current.csr[12'h3AC][31],
					ins.current.csr[12'h3AC][23],
					ins.current.csr[12'h3AC][15],
					ins.current.csr[12'h3AC][7],
					ins.current.csr[12'h3AB][31],
					ins.current.csr[12'h3AB][23],
					ins.current.csr[12'h3AB][15],
					ins.current.csr[12'h3AB][7],
					ins.current.csr[12'h3AA][31],
					ins.current.csr[12'h3AA][23],
					ins.current.csr[12'h3AA][15],
					ins.current.csr[12'h3AA][7],
					ins.current.csr[12'h3A9][31],
					ins.current.csr[12'h3A9][23],
					ins.current.csr[12'h3A9][15],
					ins.current.csr[12'h3A9][7],
					ins.current.csr[12'h3A8][31],
					ins.current.csr[12'h3A8][23],
					ins.current.csr[12'h3A8][15],
					ins.current.csr[12'h3A8][7],
					ins.current.csr[12'h3A7][31],
					ins.current.csr[12'h3A7][23],
					ins.current.csr[12'h3A7][15],
					ins.current.csr[12'h3A7][7],
					ins.current.csr[12'h3A6][31],
					ins.current.csr[12'h3A6][23],
					ins.current.csr[12'h3A6][15],
					ins.current.csr[12'h3A6][7],
					ins.current.csr[12'h3A5][31],
					ins.current.csr[12'h3A5][23],
					ins.current.csr[12'h3A5][15],
					ins.current.csr[12'h3A5][7],
					ins.current.csr[12'h3A4][31],
					ins.current.csr[12'h3A4][23],
					ins.current.csr[12'h3A4][15],
					ins.current.csr[12'h3A4][7],
					ins.current.csr[12'h3A3][31]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_L =  {
					ins.current.csr[12'h3AE][55],
					ins.current.csr[12'h3AE][47],
					ins.current.csr[12'h3AE][39],
					ins.current.csr[12'h3AE][31],
					ins.current.csr[12'h3AE][23],
					ins.current.csr[12'h3AE][15],
					ins.current.csr[12'h3AE][7],
					ins.current.csr[12'h3AC][63],
					ins.current.csr[12'h3AC][55],
					ins.current.csr[12'h3AC][47],
					ins.current.csr[12'h3AC][39],
					ins.current.csr[12'h3AC][31],
					ins.current.csr[12'h3AC][23],
					ins.current.csr[12'h3AC][15],
					ins.current.csr[12'h3AC][7],
					ins.current.csr[12'h3AA][63],
					ins.current.csr[12'h3AA][55],
					ins.current.csr[12'h3AA][47],
					ins.current.csr[12'h3AA][39],
					ins.current.csr[12'h3AA][31],
					ins.current.csr[12'h3AA][23],
					ins.current.csr[12'h3AA][15],
					ins.current.csr[12'h3AA][7],
					ins.current.csr[12'h3A8][63],
					ins.current.csr[12'h3A8][55],
					ins.current.csr[12'h3A8][47],
					ins.current.csr[12'h3A8][39],
					ins.current.csr[12'h3A8][31],
					ins.current.csr[12'h3A8][23],
					ins.current.csr[12'h3A8][15],
					ins.current.csr[12'h3A8][7],
					ins.current.csr[12'h3A6][63],
					ins.current.csr[12'h3A6][55],
					ins.current.csr[12'h3A6][47],
					ins.current.csr[12'h3A6][39],
					ins.current.csr[12'h3A6][31],
					ins.current.csr[12'h3A6][23],
					ins.current.csr[12'h3A6][15],
					ins.current.csr[12'h3A6][7],
					ins.current.csr[12'h3A4][63],
					ins.current.csr[12'h3A4][55],
					ins.current.csr[12'h3A4][47],
					ins.current.csr[12'h3A4][39],
					ins.current.csr[12'h3A4][31],
					ins.current.csr[12'h3A4][23],
					ins.current.csr[12'h3A4][15],
					ins.current.csr[12'h3A4][7],
					ins.current.csr[12'h3A2][63]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_l =  {
					ins.current.csr[12'h3A3][23],
					ins.current.csr[12'h3A3][15],
					ins.current.csr[12'h3A3][7],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A1][31],
					ins.current.csr[12'h3A1][23],
					ins.current.csr[12'h3A1][15],
					ins.current.csr[12'h3A1][7],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_l =  {
					ins.current.csr[12'h3A2][55],
					ins.current.csr[12'h3A2][47],
					ins.current.csr[12'h3A2][39],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A0][63],
					ins.current.csr[12'h3A0][55],
					ins.current.csr[12'h3A0][47],
					ins.current.csr[12'h3A0][39],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif
	PMPM_cg.sample(ins, pmpcfg, pmpaddr, pack_pmpaddr, pmpcfg_wr, pmpcfg_WR, pmpcfg_a, pmpcfg_A, pmpcfg_x, pmpcfg_X, pmpcfg_l, pmpcfg_L, pmp_hit, pmp_HIT);
endfunction
