///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_RV32PMP
covergroup RV32PMP_Baseline0_cg with function sample(ins_t ins);
    option.per_instance = 0;
    `include  "coverage/RISCV_coverage_standard_coverpoints.svh"

    read_acc: coverpoint ins.current.read_access {
        bins set = {1};
    }
    write_acc: coverpoint ins.current.write_access {
        bins set = {1};
    }
    exec_acc: coverpoint ins.current.execute_access {
        bins set = {1};
    }

    mpp_mstatus: coverpoint ins.prev.csr[12'h300][12:11] {
        bins U_mode = {2'b00};
        bins S_mode = {2'b01};
        bins M_mode = {2'b11};
    }

    Mcause:coverpoint ins.current.csr[12'h342] { 
      bins instruction_access_fault = {32'd1}; 
      bins load_access_fault        = {32'd5}; 
      bins store_access_fault       = {32'd7}; 
    }

    pmpcfg0_configurations:coverpoint ins.current.csr[12'h3A0] {
        wildcard bins no_read_pmp0cfg  = {32'b???????????????????????????????0};
        wildcard bins no_write_pmp0cfg = {32'b??????????????????????????????0?};
        wildcard bins no_exec_pmp0cfg  = {32'b?????????????????????????????0??};
        wildcard bins no_read_pmp1cfg  = {32'b???????????????????????0????????};
        wildcard bins no_write_pmp1cfg = {32'b??????????????????????0?????????};
        wildcard bins no_exec_pmp1cfg  = {32'b?????????????????????0??????????};
        wildcard bins no_read_pmp2cfg  = {32'b???????????????0????????????????};
        wildcard bins no_write_pmp2cfg = {32'b??????????????0?????????????????};
        wildcard bins no_exec_pmp2cfg  = {32'b?????????????0??????????????????};
        wildcard bins no_read_pmp3cfg  = {32'b???????0????????????????????????};
        wildcard bins no_write_pmp3cfg = {32'b??????0?????????????????????????};
        wildcard bins no_exec_pmp3cfg  = {32'b?????0??????????????????????????};
    }

    // cfg.26
    pmpcfg0_walking_ones: coverpoint ins.current.csr[12'h3A0] {
        wildcard bins walking_0  = {32'b???????????????????????????????1};
        wildcard bins walking_1  = {32'b??????????????????????????????1?};
        wildcard bins walking_2  = {32'b?????????????????????????????1??};
        wildcard bins walking_3  = {32'b????????????????????????????1???};
        wildcard bins walking_4  = {32'b???????????????????????????1????};
        wildcard bins walking_5  = {32'b??????????????????????????1?????};
        wildcard bins walking_6  = {32'b?????????????????????????1??????};
        wildcard bins walking_7  = {32'b????????????????????????1???????};
        wildcard bins walking_8  = {32'b???????????????????????1????????};
        wildcard bins walking_9  = {32'b??????????????????????1?????????};
        wildcard bins walking_10 = {32'b?????????????????????1??????????};
        wildcard bins walking_11 = {32'b????????????????????1???????????};
        wildcard bins walking_12 = {32'b???????????????????1????????????};
        wildcard bins walking_13 = {32'b??????????????????1?????????????};
        wildcard bins walking_14 = {32'b?????????????????1??????????????};
        wildcard bins walking_15 = {32'b????????????????1???????????????};
        wildcard bins walking_16 = {32'b???????????????1????????????????};
        wildcard bins walking_17 = {32'b??????????????1?????????????????};
        wildcard bins walking_18 = {32'b?????????????1??????????????????};
        wildcard bins walking_19 = {32'b????????????1???????????????????};
        wildcard bins walking_20 = {32'b???????????1????????????????????};
        wildcard bins walking_21 = {32'b??????????1?????????????????????};
        wildcard bins walking_22 = {32'b?????????1??????????????????????};
        wildcard bins walking_23 = {32'b????????1???????????????????????};
        wildcard bins walking_24 = {32'b???????1????????????????????????};
        wildcard bins walking_25 = {32'b??????1?????????????????????????};
        wildcard bins walking_26 = {32'b?????1??????????????????????????};
        wildcard bins walking_27 = {32'b????1???????????????????????????};
        wildcard bins walking_28 = {32'b???1????????????????????????????};
        wildcard bins walking_29 = {32'b??1?????????????????????????????};
        wildcard bins walking_30 = {32'b?1??????????????????????????????};
        wildcard bins walking_31 = {32'b1???????????????????????????????};        
    }

    pmpcfg0_walking_zeros: coverpoint ins.current.csr[12'h3A0] {
        wildcard bins walking_0  = {32'b???????????????????????????????0};
        wildcard bins walking_1  = {32'b??????????????????????????????0?};
        wildcard bins walking_2  = {32'b?????????????????????????????0??};
        wildcard bins walking_3  = {32'b????????????????????????????0???};
        wildcard bins walking_4  = {32'b???????????????????????????0????};
        wildcard bins walking_5  = {32'b??????????????????????????0?????};
        wildcard bins walking_6  = {32'b?????????????????????????0??????};
        wildcard bins walking_7  = {32'b????????????????????????0???????};
        wildcard bins walking_8  = {32'b???????????????????????0????????};
        wildcard bins walking_9  = {32'b??????????????????????0?????????};
        wildcard bins walking_10 = {32'b?????????????????????0??????????};
        wildcard bins walking_11 = {32'b????????????????????0???????????};
        wildcard bins walking_12 = {32'b???????????????????0????????????};
        wildcard bins walking_13 = {32'b??????????????????0?????????????};
        wildcard bins walking_14 = {32'b?????????????????0??????????????};
        wildcard bins walking_15 = {32'b????????????????0???????????????};
        wildcard bins walking_16 = {32'b???????????????0????????????????};
        wildcard bins walking_17 = {32'b??????????????0?????????????????};
        wildcard bins walking_18 = {32'b?????????????0??????????????????};
        wildcard bins walking_19 = {32'b????????????0???????????????????};
        wildcard bins walking_20 = {32'b???????????0????????????????????};
        wildcard bins walking_21 = {32'b??????????0?????????????????????};
        wildcard bins walking_22 = {32'b?????????0??????????????????????};
        wildcard bins walking_23 = {32'b????????0???????????????????????};
        wildcard bins walking_24 = {32'b???????0????????????????????????};
        wildcard bins walking_25 = {32'b??????0?????????????????????????};
        wildcard bins walking_26 = {32'b?????0??????????????????????????};
        wildcard bins walking_27 = {32'b????0???????????????????????????};
        wildcard bins walking_28 = {32'b???0????????????????????????????};
        wildcard bins walking_29 = {32'b??0?????????????????????????????};
        wildcard bins walking_30 = {32'b?0??????????????????????????????};
        wildcard bins walking_31 = {32'b0???????????????????????????????};        
    }

    // addr.3
    pmpaddr0_walking_ones: coverpoint ins.current.csr[12'h3B0] {
        wildcard bins walking_0  = {32'b???????????????????????????????1};
        wildcard bins walking_1  = {32'b??????????????????????????????1?};
        wildcard bins walking_2  = {32'b?????????????????????????????1??};
        wildcard bins walking_3  = {32'b????????????????????????????1???};
        wildcard bins walking_4  = {32'b???????????????????????????1????};
        wildcard bins walking_5  = {32'b??????????????????????????1?????};
        wildcard bins walking_6  = {32'b?????????????????????????1??????};
        wildcard bins walking_7  = {32'b????????????????????????1???????};
        wildcard bins walking_8  = {32'b???????????????????????1????????};
        wildcard bins walking_9  = {32'b??????????????????????1?????????};
        wildcard bins walking_10 = {32'b?????????????????????1??????????};
        wildcard bins walking_11 = {32'b????????????????????1???????????};
        wildcard bins walking_12 = {32'b???????????????????1????????????};
        wildcard bins walking_13 = {32'b??????????????????1?????????????};
        wildcard bins walking_14 = {32'b?????????????????1??????????????};
        wildcard bins walking_15 = {32'b????????????????1???????????????};
        wildcard bins walking_16 = {32'b???????????????1????????????????};
        wildcard bins walking_17 = {32'b??????????????1?????????????????};
        wildcard bins walking_18 = {32'b?????????????1??????????????????};
        wildcard bins walking_19 = {32'b????????????1???????????????????};
        wildcard bins walking_20 = {32'b???????????1????????????????????};
        wildcard bins walking_21 = {32'b??????????1?????????????????????};
        wildcard bins walking_22 = {32'b?????????1??????????????????????};
        wildcard bins walking_23 = {32'b????????1???????????????????????};
        wildcard bins walking_24 = {32'b???????1????????????????????????};
        wildcard bins walking_25 = {32'b??????1?????????????????????????};
        wildcard bins walking_26 = {32'b?????1??????????????????????????};
        wildcard bins walking_27 = {32'b????1???????????????????????????};
        wildcard bins walking_28 = {32'b???1????????????????????????????};
        wildcard bins walking_29 = {32'b??1?????????????????????????????};
        wildcard bins walking_30 = {32'b?1??????????????????????????????};
        wildcard bins walking_31 = {32'b1???????????????????????????????};        
    }

    pmpaddr0_walking_zeros: coverpoint ins.current.csr[12'h3B0] {
        wildcard bins walking_0  = {32'b???????????????????????????????0};
        wildcard bins walking_1  = {32'b??????????????????????????????0?};
        wildcard bins walking_2  = {32'b?????????????????????????????0??};
        wildcard bins walking_3  = {32'b????????????????????????????0???};
        wildcard bins walking_4  = {32'b???????????????????????????0????};
        wildcard bins walking_5  = {32'b??????????????????????????0?????};
        wildcard bins walking_6  = {32'b?????????????????????????0??????};
        wildcard bins walking_7  = {32'b????????????????????????0???????};
        wildcard bins walking_8  = {32'b???????????????????????0????????};
        wildcard bins walking_9  = {32'b??????????????????????0?????????};
        wildcard bins walking_10 = {32'b?????????????????????0??????????};
        wildcard bins walking_11 = {32'b????????????????????0???????????};
        wildcard bins walking_12 = {32'b???????????????????0????????????};
        wildcard bins walking_13 = {32'b??????????????????0?????????????};
        wildcard bins walking_14 = {32'b?????????????????0??????????????};
        wildcard bins walking_15 = {32'b????????????????0???????????????};
        wildcard bins walking_16 = {32'b???????????????0????????????????};
        wildcard bins walking_17 = {32'b??????????????0?????????????????};
        wildcard bins walking_18 = {32'b?????????????0??????????????????};
        wildcard bins walking_19 = {32'b????????????0???????????????????};
        wildcard bins walking_20 = {32'b???????????0????????????????????};
        wildcard bins walking_21 = {32'b??????????0?????????????????????};
        wildcard bins walking_22 = {32'b?????????0??????????????????????};
        wildcard bins walking_23 = {32'b????????0???????????????????????};
        wildcard bins walking_24 = {32'b???????0????????????????????????};
        wildcard bins walking_25 = {32'b??????0?????????????????????????};
        wildcard bins walking_26 = {32'b?????0??????????????????????????};
        wildcard bins walking_27 = {32'b????0???????????????????????????};
        wildcard bins walking_28 = {32'b???0????????????????????????????};
        wildcard bins walking_29 = {32'b??0?????????????????????????????};
        wildcard bins walking_30 = {32'b?0??????????????????????????????};
        wildcard bins walking_31 = {32'b0???????????????????????????????};        
    }

    pmpaddr1_walking_ones: coverpoint ins.current.csr[12'h3B1] {
        wildcard bins walking_0  = {32'b???????????????????????????????1};
        wildcard bins walking_1  = {32'b??????????????????????????????1?};
        wildcard bins walking_2  = {32'b?????????????????????????????1??};
        wildcard bins walking_3  = {32'b????????????????????????????1???};
        wildcard bins walking_4  = {32'b???????????????????????????1????};
        wildcard bins walking_5  = {32'b??????????????????????????1?????};
        wildcard bins walking_6  = {32'b?????????????????????????1??????};
        wildcard bins walking_7  = {32'b????????????????????????1???????};
        wildcard bins walking_8  = {32'b???????????????????????1????????};
        wildcard bins walking_9  = {32'b??????????????????????1?????????};
        wildcard bins walking_10 = {32'b?????????????????????1??????????};
        wildcard bins walking_11 = {32'b????????????????????1???????????};
        wildcard bins walking_12 = {32'b???????????????????1????????????};
        wildcard bins walking_13 = {32'b??????????????????1?????????????};
        wildcard bins walking_14 = {32'b?????????????????1??????????????};
        wildcard bins walking_15 = {32'b????????????????1???????????????};
        wildcard bins walking_16 = {32'b???????????????1????????????????};
        wildcard bins walking_17 = {32'b??????????????1?????????????????};
        wildcard bins walking_18 = {32'b?????????????1??????????????????};
        wildcard bins walking_19 = {32'b????????????1???????????????????};
        wildcard bins walking_20 = {32'b???????????1????????????????????};
        wildcard bins walking_21 = {32'b??????????1?????????????????????};
        wildcard bins walking_22 = {32'b?????????1??????????????????????};
        wildcard bins walking_23 = {32'b????????1???????????????????????};
        wildcard bins walking_24 = {32'b???????1????????????????????????};
        wildcard bins walking_25 = {32'b??????1?????????????????????????};
        wildcard bins walking_26 = {32'b?????1??????????????????????????};
        wildcard bins walking_27 = {32'b????1???????????????????????????};
        wildcard bins walking_28 = {32'b???1????????????????????????????};
        wildcard bins walking_29 = {32'b??1?????????????????????????????};
        wildcard bins walking_30 = {32'b?1??????????????????????????????};
        wildcard bins walking_31 = {32'b1???????????????????????????????};        
    }

    pmpaddr1_walking_zeros: coverpoint ins.current.csr[12'h3B1] {
        wildcard bins walking_0  = {32'b???????????????????????????????0};
        wildcard bins walking_1  = {32'b??????????????????????????????0?};
        wildcard bins walking_2  = {32'b?????????????????????????????0??};
        wildcard bins walking_3  = {32'b????????????????????????????0???};
        wildcard bins walking_4  = {32'b???????????????????????????0????};
        wildcard bins walking_5  = {32'b??????????????????????????0?????};
        wildcard bins walking_6  = {32'b?????????????????????????0??????};
        wildcard bins walking_7  = {32'b????????????????????????0???????};
        wildcard bins walking_8  = {32'b???????????????????????0????????};
        wildcard bins walking_9  = {32'b??????????????????????0?????????};
        wildcard bins walking_10 = {32'b?????????????????????0??????????};
        wildcard bins walking_11 = {32'b????????????????????0???????????};
        wildcard bins walking_12 = {32'b???????????????????0????????????};
        wildcard bins walking_13 = {32'b??????????????????0?????????????};
        wildcard bins walking_14 = {32'b?????????????????0??????????????};
        wildcard bins walking_15 = {32'b????????????????0???????????????};
        wildcard bins walking_16 = {32'b???????????????0????????????????};
        wildcard bins walking_17 = {32'b??????????????0?????????????????};
        wildcard bins walking_18 = {32'b?????????????0??????????????????};
        wildcard bins walking_19 = {32'b????????????0???????????????????};
        wildcard bins walking_20 = {32'b???????????0????????????????????};
        wildcard bins walking_21 = {32'b??????????0?????????????????????};
        wildcard bins walking_22 = {32'b?????????0??????????????????????};
        wildcard bins walking_23 = {32'b????????0???????????????????????};
        wildcard bins walking_24 = {32'b???????0????????????????????????};
        wildcard bins walking_25 = {32'b??????0?????????????????????????};
        wildcard bins walking_26 = {32'b?????0??????????????????????????};
        wildcard bins walking_27 = {32'b????0???????????????????????????};
        wildcard bins walking_28 = {32'b???0????????????????????????????};
        wildcard bins walking_29 = {32'b??0?????????????????????????????};
        wildcard bins walking_30 = {32'b?0??????????????????????????????};
        wildcard bins walking_31 = {32'b0???????????????????????????????};        
    }

    pmpaddr2_walking_ones: coverpoint ins.current.csr[12'h3B2] {
        wildcard bins walking_0  = {32'b???????????????????????????????1};
        wildcard bins walking_1  = {32'b??????????????????????????????1?};
        wildcard bins walking_2  = {32'b?????????????????????????????1??};
        wildcard bins walking_3  = {32'b????????????????????????????1???};
        wildcard bins walking_4  = {32'b???????????????????????????1????};
        wildcard bins walking_5  = {32'b??????????????????????????1?????};
        wildcard bins walking_6  = {32'b?????????????????????????1??????};
        wildcard bins walking_7  = {32'b????????????????????????1???????};
        wildcard bins walking_8  = {32'b???????????????????????1????????};
        wildcard bins walking_9  = {32'b??????????????????????1?????????};
        wildcard bins walking_10 = {32'b?????????????????????1??????????};
        wildcard bins walking_11 = {32'b????????????????????1???????????};
        wildcard bins walking_12 = {32'b???????????????????1????????????};
        wildcard bins walking_13 = {32'b??????????????????1?????????????};
        wildcard bins walking_14 = {32'b?????????????????1??????????????};
        wildcard bins walking_15 = {32'b????????????????1???????????????};
        wildcard bins walking_16 = {32'b???????????????1????????????????};
        wildcard bins walking_17 = {32'b??????????????1?????????????????};
        wildcard bins walking_18 = {32'b?????????????1??????????????????};
        wildcard bins walking_19 = {32'b????????????1???????????????????};
        wildcard bins walking_20 = {32'b???????????1????????????????????};
        wildcard bins walking_21 = {32'b??????????1?????????????????????};
        wildcard bins walking_22 = {32'b?????????1??????????????????????};
        wildcard bins walking_23 = {32'b????????1???????????????????????};
        wildcard bins walking_24 = {32'b???????1????????????????????????};
        wildcard bins walking_25 = {32'b??????1?????????????????????????};
        wildcard bins walking_26 = {32'b?????1??????????????????????????};
        wildcard bins walking_27 = {32'b????1???????????????????????????};
        wildcard bins walking_28 = {32'b???1????????????????????????????};
        wildcard bins walking_29 = {32'b??1?????????????????????????????};
        wildcard bins walking_30 = {32'b?1??????????????????????????????};
        wildcard bins walking_31 = {32'b1???????????????????????????????};        
    }

    pmpaddr2_walking_zeros: coverpoint ins.current.csr[12'h3B2] {
        wildcard bins walking_0  = {32'b???????????????????????????????0};
        wildcard bins walking_1  = {32'b??????????????????????????????0?};
        wildcard bins walking_2  = {32'b?????????????????????????????0??};
        wildcard bins walking_3  = {32'b????????????????????????????0???};
        wildcard bins walking_4  = {32'b???????????????????????????0????};
        wildcard bins walking_5  = {32'b??????????????????????????0?????};
        wildcard bins walking_6  = {32'b?????????????????????????0??????};
        wildcard bins walking_7  = {32'b????????????????????????0???????};
        wildcard bins walking_8  = {32'b???????????????????????0????????};
        wildcard bins walking_9  = {32'b??????????????????????0?????????};
        wildcard bins walking_10 = {32'b?????????????????????0??????????};
        wildcard bins walking_11 = {32'b????????????????????0???????????};
        wildcard bins walking_12 = {32'b???????????????????0????????????};
        wildcard bins walking_13 = {32'b??????????????????0?????????????};
        wildcard bins walking_14 = {32'b?????????????????0??????????????};
        wildcard bins walking_15 = {32'b????????????????0???????????????};
        wildcard bins walking_16 = {32'b???????????????0????????????????};
        wildcard bins walking_17 = {32'b??????????????0?????????????????};
        wildcard bins walking_18 = {32'b?????????????0??????????????????};
        wildcard bins walking_19 = {32'b????????????0???????????????????};
        wildcard bins walking_20 = {32'b???????????0????????????????????};
        wildcard bins walking_21 = {32'b??????????0?????????????????????};
        wildcard bins walking_22 = {32'b?????????0??????????????????????};
        wildcard bins walking_23 = {32'b????????0???????????????????????};
        wildcard bins walking_24 = {32'b???????0????????????????????????};
        wildcard bins walking_25 = {32'b??????0?????????????????????????};
        wildcard bins walking_26 = {32'b?????0??????????????????????????};
        wildcard bins walking_27 = {32'b????0???????????????????????????};
        wildcard bins walking_28 = {32'b???0????????????????????????????};
        wildcard bins walking_29 = {32'b??0?????????????????????????????};
        wildcard bins walking_30 = {32'b?0??????????????????????????????};
        wildcard bins walking_31 = {32'b0???????????????????????????????};        
    }

    pmpaddr3_walking_ones: coverpoint ins.current.csr[12'h3B3] {
        wildcard bins walking_0  = {32'b???????????????????????????????1};
        wildcard bins walking_1  = {32'b??????????????????????????????1?};
        wildcard bins walking_2  = {32'b?????????????????????????????1??};
        wildcard bins walking_3  = {32'b????????????????????????????1???};
        wildcard bins walking_4  = {32'b???????????????????????????1????};
        wildcard bins walking_5  = {32'b??????????????????????????1?????};
        wildcard bins walking_6  = {32'b?????????????????????????1??????};
        wildcard bins walking_7  = {32'b????????????????????????1???????};
        wildcard bins walking_8  = {32'b???????????????????????1????????};
        wildcard bins walking_9  = {32'b??????????????????????1?????????};
        wildcard bins walking_10 = {32'b?????????????????????1??????????};
        wildcard bins walking_11 = {32'b????????????????????1???????????};
        wildcard bins walking_12 = {32'b???????????????????1????????????};
        wildcard bins walking_13 = {32'b??????????????????1?????????????};
        wildcard bins walking_14 = {32'b?????????????????1??????????????};
        wildcard bins walking_15 = {32'b????????????????1???????????????};
        wildcard bins walking_16 = {32'b???????????????1????????????????};
        wildcard bins walking_17 = {32'b??????????????1?????????????????};
        wildcard bins walking_18 = {32'b?????????????1??????????????????};
        wildcard bins walking_19 = {32'b????????????1???????????????????};
        wildcard bins walking_20 = {32'b???????????1????????????????????};
        wildcard bins walking_21 = {32'b??????????1?????????????????????};
        wildcard bins walking_22 = {32'b?????????1??????????????????????};
        wildcard bins walking_23 = {32'b????????1???????????????????????};
        wildcard bins walking_24 = {32'b???????1????????????????????????};
        wildcard bins walking_25 = {32'b??????1?????????????????????????};
        wildcard bins walking_26 = {32'b?????1??????????????????????????};
        wildcard bins walking_27 = {32'b????1???????????????????????????};
        wildcard bins walking_28 = {32'b???1????????????????????????????};
        wildcard bins walking_29 = {32'b??1?????????????????????????????};
        wildcard bins walking_30 = {32'b?1??????????????????????????????};
        wildcard bins walking_31 = {32'b1???????????????????????????????};        
    }

    pmpaddr3_walking_zeros: coverpoint ins.current.csr[12'h3B3] {
        wildcard bins walking_0  = {32'b???????????????????????????????0};
        wildcard bins walking_1  = {32'b??????????????????????????????0?};
        wildcard bins walking_2  = {32'b?????????????????????????????0??};
        wildcard bins walking_3  = {32'b????????????????????????????0???};
        wildcard bins walking_4  = {32'b???????????????????????????0????};
        wildcard bins walking_5  = {32'b??????????????????????????0?????};
        wildcard bins walking_6  = {32'b?????????????????????????0??????};
        wildcard bins walking_7  = {32'b????????????????????????0???????};
        wildcard bins walking_8  = {32'b???????????????????????0????????};
        wildcard bins walking_9  = {32'b??????????????????????0?????????};
        wildcard bins walking_10 = {32'b?????????????????????0??????????};
        wildcard bins walking_11 = {32'b????????????????????0???????????};
        wildcard bins walking_12 = {32'b???????????????????0????????????};
        wildcard bins walking_13 = {32'b??????????????????0?????????????};
        wildcard bins walking_14 = {32'b?????????????????0??????????????};
        wildcard bins walking_15 = {32'b????????????????0???????????????};
        wildcard bins walking_16 = {32'b???????????????0????????????????};
        wildcard bins walking_17 = {32'b??????????????0?????????????????};
        wildcard bins walking_18 = {32'b?????????????0??????????????????};
        wildcard bins walking_19 = {32'b????????????0???????????????????};
        wildcard bins walking_20 = {32'b???????????0????????????????????};
        wildcard bins walking_21 = {32'b??????????0?????????????????????};
        wildcard bins walking_22 = {32'b?????????0??????????????????????};
        wildcard bins walking_23 = {32'b????????0???????????????????????};
        wildcard bins walking_24 = {32'b???????0????????????????????????};
        wildcard bins walking_25 = {32'b??????0?????????????????????????};
        wildcard bins walking_26 = {32'b?????0??????????????????????????};
        wildcard bins walking_27 = {32'b????0???????????????????????????};
        wildcard bins walking_28 = {32'b???0????????????????????????????};
        wildcard bins walking_29 = {32'b??0?????????????????????????????};
        wildcard bins walking_30 = {32'b?0??????????????????????????????};
        wildcard bins walking_31 = {32'b0???????????????????????????????};        
    }

    instr_acc_fault: cross mpp_mstatus, exec_acc, pmpcfg0_configurations, Mcause { // exp.1
        ignore_bins ig1  = binsof(Mcause.load_access_fault);
        ignore_bins ig2  = binsof(Mcause.store_access_fault);
        ignore_bins ig3  = binsof(pmpcfg0_configurations.no_read_pmp0cfg);
        ignore_bins ig4  = binsof(pmpcfg0_configurations.no_read_pmp1cfg);
        ignore_bins ig5  = binsof(pmpcfg0_configurations.no_read_pmp2cfg);
        ignore_bins ig6  = binsof(pmpcfg0_configurations.no_read_pmp3cfg);
        ignore_bins ig7  = binsof(pmpcfg0_configurations.no_write_pmp0cfg);
        ignore_bins ig8  = binsof(pmpcfg0_configurations.no_write_pmp1cfg);
        ignore_bins ig9  = binsof(pmpcfg0_configurations.no_write_pmp2cfg);
        ignore_bins ig10 = binsof(pmpcfg0_configurations.no_write_pmp3cfg);
    } 

    load_acc_fault: cross mpp_mstatus, read_acc, pmpcfg0_configurations, Mcause { // exp.2
        ignore_bins ig1 = binsof(Mcause.instruction_access_fault);
        ignore_bins ig2 = binsof(Mcause.store_access_fault);
        ignore_bins ig3  = binsof(pmpcfg0_configurations.no_exec_pmp0cfg);
        ignore_bins ig4  = binsof(pmpcfg0_configurations.no_exec_pmp1cfg);
        ignore_bins ig5  = binsof(pmpcfg0_configurations.no_exec_pmp2cfg);
        ignore_bins ig6  = binsof(pmpcfg0_configurations.no_exec_pmp3cfg);
        ignore_bins ig7  = binsof(pmpcfg0_configurations.no_write_pmp0cfg);
        ignore_bins ig8  = binsof(pmpcfg0_configurations.no_write_pmp1cfg);
        ignore_bins ig9  = binsof(pmpcfg0_configurations.no_write_pmp2cfg);
        ignore_bins ig10 = binsof(pmpcfg0_configurations.no_write_pmp3cfg);
    }

    store_acc_fault: cross mpp_mstatus, write_acc, pmpcfg0_configurations, Mcause { // exp.3
        ignore_bins ig1 = binsof(Mcause.instruction_access_fault);
        ignore_bins ig2 = binsof(Mcause.load_access_fault);
        ignore_bins ig3  = binsof(pmpcfg0_configurations.no_read_pmp0cfg);
        ignore_bins ig4  = binsof(pmpcfg0_configurations.no_read_pmp1cfg);
        ignore_bins ig5  = binsof(pmpcfg0_configurations.no_read_pmp2cfg);
        ignore_bins ig6  = binsof(pmpcfg0_configurations.no_read_pmp3cfg);
        ignore_bins ig7  = binsof(pmpcfg0_configurations.no_exec_pmp0cfg);
        ignore_bins ig8  = binsof(pmpcfg0_configurations.no_exec_pmp1cfg);
        ignore_bins ig9  = binsof(pmpcfg0_configurations.no_exec_pmp2cfg);
        ignore_bins ig10 = binsof(pmpcfg0_configurations.no_exec_pmp3cfg);
    }
endgroup

function void rv32pmp_sample(int hart, int issue, ins_t ins);
    RV32PMP_Baseline0_cg.sample(ins);
endfunction
