///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    c_lbu_cg = new(); c_lbu_cg.set_inst_name("obj_c_lbu");
    c_lh_cg = new(); c_lh_cg.set_inst_name("obj_c_lh");
    c_lhu_cg = new(); c_lhu_cg.set_inst_name("obj_c_lhu");
    c_not_cg = new(); c_not_cg.set_inst_name("obj_c_not");
    c_sb_cg = new(); c_sb_cg.set_inst_name("obj_c_sb");
    c_sh_cg = new(); c_sh_cg.set_inst_name("obj_c_sh");
    c_zext_b_cg = new(); c_zext_b_cg.set_inst_name("obj_c_zext_b");
