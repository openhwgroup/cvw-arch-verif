///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_RV64ZCBZBB
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_rv64zcbzbb_t;


covergroup c_sext_b_cg with function sample(ins_rv64zcbzbb_t ins);
    option.per_instance = 1; 
    option.comment = "c.sext.b";
    cp_asm_count : coverpoint ins.ins_str == "sext.b"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rdp : coverpoint ins.get_gpr_c_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rd_corners_lb : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111111111111111111111111111110000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111111111111111111111111111110000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000000000001111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000000000001111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111111111111111111111111111110101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000000000000000000000000000001010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000000000001011011};
        wildcard bins random1  = {64'b1111111111111111111111111111111111111111111111111111111111011011}; 
     }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1p : coverpoint ins.get_gpr_c_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
endgroup

covergroup c_sext_h_cg with function sample(ins_rv64zcbzbb_t ins);
    option.per_instance = 1; 
    option.comment = "c.sext.h";
    cp_asm_count : coverpoint ins.ins_str == "sext.h"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rdp : coverpoint ins.get_gpr_c_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
cp_rd_corners_lh : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111111111111111111111000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111111111111111111111000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b0000000000000000000000000000000000000000000000000101010101010101};
        wildcard bins walkeven = {64'b1111111111111111111111111111111111111111111111111010101010101010};
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000101101110111100};
        wildcard bins random1  = {64'b1111111111111111111111111111111111111111111111111101101110111100};
     }    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1p : coverpoint ins.get_gpr_c_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
endgroup

covergroup c_zext_h_cg with function sample(ins_rv64zcbzbb_t ins);
    option.per_instance = 1; 
    option.comment = "c.zext.h";
    cp_asm_count : coverpoint ins.ins_str == "zext.h"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rdp : coverpoint ins.get_gpr_c_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
cp_rd_corners_lhu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0)  {
        option.comment = "RD Corners";
        wildcard bins zero     = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b0000000000000000000000000000000000000000000000001000000000000000};        // Zero Extended min half word
        wildcard bins minp1    = {64'b0000000000000000000000000000000000000000000000001000000000000001};        // Zero Extended minp1 half word
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000111111111111111};        // Zero Extended max half word
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000111111111111110};        // Zero Extended maxm1 half word
        wildcard bins ones     = {64'b0000000000000000000000000000000000000000000000001111111111111111};        // Zero Extended ones half word
        wildcard bins onesm1   = {64'b0000000000000000000000000000000000000000000000001111111111111110};        // Zero Extended onesm1 half word
        wildcard bins walkeodd = {64'b0000000000000000000000000000000000000000000000000101010101010101};        // Zero Extended walkodd
        wildcard bins walkeven = {64'b0000000000000000000000000000000000000000000000001010101010101010};        // Zero Extended walkeven
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000101101110111100};        // Zero Extended random1
        wildcard bins random1  = {64'b0000000000000000000000000000000000000000000000001101101110111100};        // Zero Extended random1
     }    cp_rd_toggle_lhu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
    }
    cp_rs1p : coverpoint ins.get_gpr_c_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
endgroup

function void rv64zcbzbb_sample(int hart, int issue);
    ins_rv64zcbzbb_t ins;
    if (traceDataQ[hart][issue][0].insn[1:0] != 3) begin // compressed instruction
        $display("Examining compressed instruction rv64zcbzbb_sample with inst_name = %s disass = %s", traceDataQ[hart][issue][0].inst_name, traceDataQ[hart][issue][0].disass);
        case (traceDataQ[hart][issue][0].inst_name)
            "sext.b" : begin
                if (traceDataQ[hart][issue][0].insn[1:0] == 2'b01 && traceDataQ[hart][issue][0].insn[6:2] == 5'b11001) begin // Specific bits for "sext.b"
                    ins = new(hart, issue, traceDataQ);
                    ins.add_rd(0);      
                    ins.add_rs1(1);     
                    c_sext_b_cg.sample(ins); 
                end
            end
            "zext.h" : begin
                if (traceDataQ[hart][issue][0].insn[1:0] == 2'b01 && traceDataQ[hart][issue][0].insn[6:2] == 5'b11010) begin // Specific bits for "zext.h"
                    ins = new(hart, issue, traceDataQ);
                    ins.add_rd(0);       
                    ins.add_rs1(1);     
                    c_zext_h_cg.sample(ins); 
                end
            end
            "sext.h" : begin
                if (traceDataQ[hart][issue][0].insn[1:0] == 2'b01 && traceDataQ[hart][issue][0].insn[6:2] == 5'b11011) begin // Specific bits for "sext.h"
                    ins = new(hart, issue, traceDataQ);
                    ins.add_rd(0);       
                    ins.add_rs1(1);      
                    c_sext_h_cg.sample(ins); 
                end
            end
        endcase
    end
endfunction
