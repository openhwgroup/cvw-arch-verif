///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fcsr_cg = new();         fcsr_cg.set_inst_name("obj_fcsr");
    frm_cg = new();         frm_cg.set_inst_name("obj_frm");
    fflags_cg = new();       fflags_cg.set_inst_name("obj_fflags");
