///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    c_flw_cg = new(); c_flw_cg.set_inst_name("obj_c_flw");
    c_flwsp_cg = new(); c_flwsp_cg.set_inst_name("obj_c_flwsp");
    c_fsw_cg = new(); c_fsw_cg.set_inst_name("obj_c_fsw");
    c_fswsp_cg = new(); c_fswsp_cg.set_inst_name("obj_c_fswsp");
