///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fcvt_d_h_cg = new(); fcvt_d_h_cg.set_inst_name("obj_fcvt_d_h");
    fcvt_h_d_cg = new(); fcvt_h_d_cg.set_inst_name("obj_fcvt_h_d");
