///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    mcsr_cg = new();        mcsr_cg.set_inst_name("obj_mcsr");
    mcause_cg = new();      mcause_cg.set_inst_name("obj_mcause");
    mstatus_cg = new();     mstatus_cg.set_inst_name("obj_mstatus");
    mprivinst_cg = new();   mprivinst_cg.set_inst_name("obj_mprivinst");

 
