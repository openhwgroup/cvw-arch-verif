///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Written: Corey Hickson chickson@hmc.edu 23 November 2024
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_EXCEPTIONSF
covergroup ExceptionsF_exceptions_cg with function sample(ins_t ins);
    option.per_instance = 0; 

    // building blocks for the main coverpoints
    mstatus_FS_zero: coverpoint ins.prev.csr[12'h300][14:13] {
        bins disabled = {2'b00};
    }
    mstatus_FS_nonzero: coverpoint ins.prev.csr[12'h300][14:13] {
        bins enabled = {!2'b00};
    }
    frm_illegal: coverpoint ins.prev.csr[12'h003][7:5] {
        bins reserved_5 = {3'b101};
        bins reserved_6 = {3'b110};
        bins reserved_7 = {3'b111};
    }
    // csrrw: coverpoint ins.current.insn {
    //     wildcard bins csrrw = {32'b????????????_?????_001_?????_1110011}; 
    // }
    // fp_csrs: coverpoint ins.current.insn[31:20] {
    //     bins fcsr   = {12'h003};
    //     bins frm    = {12'h002};
    //     bins fflags = {12'h001};
    // }
    instrs: coverpoint ins.current.insn {
        wildcard bins fsw          = {32'b????????????_?????_010_?????_0100111};
        wildcard bins flw          = {32'b????????????_?????_010_?????_0000111};
        wildcard bins fadd         = {32'b00000_??_?????_?????_???_?????_1010011};
        wildcard bins fsub         = {32'b00001_??_?????_?????_???_?????_1010011};
        wildcard bins fmul         = {32'b00010_??_?????_?????_???_?????_1010011};
        wildcard bins fdiv         = {32'b00011_??_?????_?????_???_?????_1010011};
        wildcard bins fcvt_x_f     = {32'b11000_??_?????_?????_???_?????_1010011};
        wildcard bins fcvt_f_x     = {32'b11010_??_?????_?????_???_?????_1010011};
        wildcard bins fcvt_f_f     = {32'b01000_??_?????_?????_???_?????_1010011};
        wildcard bins fmadd        = {32'b?????_??_?????_?????_???_?????_1000011};
        wildcard bins fsqrt        = {32'b01011_??_00000_?????_???_?????_1010011};
        wildcard bins fsgnj        = {32'b00100_??_?????_?????_000_?????_1010011};
        wildcard bins feq          = {32'b10100_??_?????_?????_010_?????_1010011};
        wildcard bins fmv_x_f      = {32'b11100_??_00000_?????_000_?????_1010011};
        wildcard bins fmv_f_x      = {32'b11110_??_00000_?????_000_?????_1010011};
        wildcard bins fclass       = {32'b11100_??_00000_?????_001_?????_1010011};
        wildcard bins fmin         = {32'b00101_??_?????_?????_000_?????_1010011};
        wildcard bins fli          = {32'b11110_??_00001_?????_000_?????_1010011};
        wildcard bins fround       = {32'b01000_??_00100_?????_???_?????_1010011};
        wildcard bins add          = {32'b0000000_?????_?????_000_?????_0110011};
        wildcard bins csrrw_fcsr   = {32'b000000000011_?????_001_?????_1110011};
        wildcard bins csrrw_frm    = {32'b000000000010_?????_001_?????_1110011};
        wildcard bins csrrw_fflags = {32'b000000000001_?????_001_?????_1110011};
        wildcard bins csrrs_fcsr   = {32'b000000000011_?????_010_?????_1110011};
        wildcard bins csrrs_frm    = {32'b000000000010_?????_010_?????_1110011};
        wildcard bins csrrs_fflags = {32'b000000000001_?????_010_?????_1110011};
        wildcard bins csrrc_fcsr   = {32'b000000000011_?????_011_?????_1110011};
        wildcard bins csrrc_frm    = {32'b000000000010_?????_011_?????_1110011};
        wildcard bins csrrc_fflags = {32'b000000000001_?????_011_?????_1110011};
        `ifdef XLEN32
            wildcard bins fmvh         = {32'b1110001_00001_?????_000_?????_1010011};
            wildcard bins fmvp         = {32'b1011001_?????_?????_000_?????_1010011};
        `endif
    }
    dyn_instrs: coverpoint ins.current.insn {
        wildcard bins fadd_dyn     = {32'b00000_??_?????_?????_111_?????_1010011};
        wildcard bins fsub_dyn     = {32'b00001_??_?????_?????_111_?????_1010011};
        wildcard bins fmul_dyn     = {32'b00010_??_?????_?????_111_?????_1010011};
        wildcard bins fdiv_dyn     = {32'b00011_??_?????_?????_111_?????_1010011};
        wildcard bins fcvt_x_f_dyn = {32'b11000_??_?????_?????_111_?????_1010011};
        wildcard bins fcvt_f_f_dyn = {32'b01000_??_?????_?????_111_?????_1010011};
        wildcard bins fmadd_dyn    = {32'b?????_??_?????_?????_111_?????_1000011};
        wildcard bins fsqrt_dyn    = {32'b01011_??_00000_?????_111_?????_1010011};
        wildcard bins fround_dyn   = {32'b01000_??_00100_?????_111_?????_1010011};
    }
    // main coverpoints
    cp_mstatus_fs_illegal_instr: cross instrs, mstatus_FS_zero;
    // cp_mstatus_fs_csr_write:  redundant, covered by cp_mstatus_fs_illegal_instr
    cp_badfrm: cross dyn_instrs, mstatus_FS_nonzero, frm_illegal;
endgroup

function void exceptionsf_sample(int hart, int issue, ins_t ins);
    ExceptionsF_exceptions_cg.sample(ins);
endfunction
