///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    c_fld_cg = new(); c_fld_cg.set_inst_name("obj_c_fld");
    c_fldsp_cg = new(); c_fldsp_cg.set_inst_name("obj_c_fldsp");
    c_fsd_cg = new(); c_fsd_cg.set_inst_name("obj_c_fsd");
    c_fsdsp_cg = new(); c_fsdsp_cg.set_inst_name("obj_c_fsdsp");
