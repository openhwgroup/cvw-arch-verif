///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////
    ExceptionsV_vadd_vv_cg = new(); ExceptionsV_vadd_vv_cg.set_inst_name("obj_ExceptionsV_vadd_vv");
