///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    c_add_cg = new(); c_add_cg.set_inst_name("obj_c_add");
    c_addi_cg = new(); c_addi_cg.set_inst_name("obj_c_addi");
    c_addi16sp_cg = new(); c_addi16sp_cg.set_inst_name("obj_c_addi16sp");
    c_addi4spn_cg = new(); c_addi4spn_cg.set_inst_name("obj_c_addi4spn");
    c_addiw_cg = new(); c_addiw_cg.set_inst_name("obj_c_addiw");
    c_addw_cg = new(); c_addw_cg.set_inst_name("obj_c_addw");
    c_and_cg = new(); c_and_cg.set_inst_name("obj_c_and");
    c_andi_cg = new(); c_andi_cg.set_inst_name("obj_c_andi");
    c_beqz_cg = new(); c_beqz_cg.set_inst_name("obj_c_beqz");
    c_bnez_cg = new(); c_bnez_cg.set_inst_name("obj_c_bnez");
    c_j_cg = new(); c_j_cg.set_inst_name("obj_c_j");
    c_jalr_cg = new(); c_jalr_cg.set_inst_name("obj_c_jalr");
    c_jr_cg = new(); c_jr_cg.set_inst_name("obj_c_jr");
    c_ld_cg = new(); c_ld_cg.set_inst_name("obj_c_ld");
    c_ldsp_cg = new(); c_ldsp_cg.set_inst_name("obj_c_ldsp");
    c_li_cg = new(); c_li_cg.set_inst_name("obj_c_li");
    c_lui_cg = new(); c_lui_cg.set_inst_name("obj_c_lui");
    c_lw_cg = new(); c_lw_cg.set_inst_name("obj_c_lw");
    c_lwsp_cg = new(); c_lwsp_cg.set_inst_name("obj_c_lwsp");
    c_mv_cg = new(); c_mv_cg.set_inst_name("obj_c_mv");
    c_nop_cg = new(); c_nop_cg.set_inst_name("obj_c_nop");
    c_or_cg = new(); c_or_cg.set_inst_name("obj_c_or");
    c_sd_cg = new(); c_sd_cg.set_inst_name("obj_c_sd");
    c_sdsp_cg = new(); c_sdsp_cg.set_inst_name("obj_c_sdsp");
    c_slli_cg = new(); c_slli_cg.set_inst_name("obj_c_slli");
    c_srai_cg = new(); c_srai_cg.set_inst_name("obj_c_srai");
    c_srli_cg = new(); c_srli_cg.set_inst_name("obj_c_srli");
    c_sub_cg = new(); c_sub_cg.set_inst_name("obj_c_sub");
    c_subw_cg = new(); c_subw_cg.set_inst_name("obj_c_subw");
    c_sw_cg = new(); c_sw_cg.set_inst_name("obj_c_sw");
    c_swsp_cg = new(); c_swsp_cg.set_inst_name("obj_c_swsp");
    c_xor_cg = new(); c_xor_cg.set_inst_name("obj_c_xor");
