///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    RV64VMZicbom_cbo_inval_cg = new(); RV64VMZicbom_cbo_inval_cg.set_inst_name("obj_RV64VMZicbom_cbo_inval");
    RV64VMZicbom_cbo_clean_cg = new(); RV64VMZicbom_cbo_clean_cg.set_inst_name("obj_RV64VMZicbom_cbo_clean");
    RV64VMZicbom_cbo_flush_cg = new(); RV64VMZicbom_cbo_flush_cg.set_inst_name("obj_RV64VMZicbom_cbo_flush");