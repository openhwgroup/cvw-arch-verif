///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Standard Covergroups
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file
// except in compliance with the License, or, at your option, the Apache License version 2.0. You
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied. See the License for the specific language governing permissions
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

//------------ Assuming it right for time being --------------

`define RAMBASEADDR 32'h80000000
`define LARGESTPROGRAM 32'h00010000
`define SAFEREGIONSTART (`RAMBASEADDR + `LARGESTPROGRAM)
`define REGIONSTART `SAFEREGIONSTART

`define G 2              // Set G as needed (0, 1, 2, etc.)
`define g (2**(`G+2))    // Region size = 2^(G+2)

// Define PMP_16 or PMP_64
`define PMP_16

// --- STANDARD_REGION macro based on G value ---

// Case: G == 0    NA4 granularity (shift by 2)
`define REGION_G0    (`REGIONSTART >> 2)

// Case: G == 1    region has one trailing 0
`define STANDARD_REGION_G1    (`REGIONSTART >> (`G+2))

// Case: G >= 2    region has (G-1) trailing 1s
`define STANDARD_REGION_GX    (`REGIONSTART >> (`G+2)) | ((1 << (`G-1)) - 1)

// Alias one of the above depending on G
`define STANDARD_REGION `STANDARD_REGION_GX

//------------------------------------------------------------

`define COVER_RV32PMP
`define COVER_RV64PMP

covergroup PMPM_cg with function sample(ins_t ins, logic [XLEN-1:0] pmpcfg [15:0], logic [XLEN-1:0] pmpaddr [62:0], logic [29:0] pmpcfg_rw, logic [95:0] pmpcfg_RW, logic [29:0] pmpcfg_a, logic [95:0] pmpcfg_A, logic [14:0] pmpcfg_x, logic [47:0] pmpcfg_X, logic [14:0] pmpcfg_l, logic [47:0] pmpcfg_L, logic [14:0] pmp_hit, logic [47:0] pmp_HIT);
	option.per_instance = 0;
	`include  "coverage/RISCV_coverage_standard_coverpoints.svh"

	addr_in_region: coverpoint (ins.current.rs1_val + ins.current.imm) {
		bins at_region = {`STANDARD_REGION};
	}

	addr_offset: coverpoint (ins.current.rs1_val + ins.current.imm) {
  		bins at_base      = {`REGIONSTART};

  		// this should fault, since it’s outside the region
  		bins below_base   = {`REGIONSTART-4};

		//just into the region
  		bins above_base   = {`REGIONSTART+4};

  		// this should also fault as “outside”, but loads beyond this should succeed
  		bins just_beyond  = {`REGIONSTART+`g};

		//last word inside region
		bins highest_word  = {`REGIONSTART +`g-4};
	}

	exec_instr: coverpoint ins.current.insn {
		wildcard bins jalr = {32'b????????????_?????_000_?????_1100111};
	}

	read_instr_lw: coverpoint ins.current.insn {
		wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
	}

	read_instr: coverpoint ins.current.insn {
		wildcard bins lb  = {32'b????????????_?????_000_?????_0000011};
		wildcard bins lbu = {32'b????????????_?????_100_?????_0000011};
		wildcard bins lh  = {32'b????????????_?????_001_?????_0000011};
		wildcard bins lhu = {32'b????????????_?????_101_?????_0000011};
		wildcard bins lw  = {32'b????????????_?????_010_?????_0000011};
		`ifdef XLEN64
			wildcard bins lwu = {32'b????????????_?????_110_?????_0000011};
			wildcard bins ld  = {32'b????????????_?????_011_?????_0000011};
		`endif
	}

	write_instr_sw: coverpoint ins.current.insn {
		wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
	}

	write_instr: coverpoint ins.current.insn {
		wildcard bins sb = {32'b???????_?????_?????_000_?????_0100011};
		wildcard bins sh = {32'b???????_?????_?????_001_?????_0100011};
		wildcard bins sw = {32'b???????_?????_?????_010_?????_0100011};
		`ifdef XLEN64
			wildcard bins sd = {32'b???????_?????_?????_011_?????_0100011};
		`endif
	}

//-------------------------------------------------------

	standard_region: coverpoint pmpaddr[0] {
		bins standard_region = {`STANDARD_REGION};
	}

	legal_lxwr: coverpoint pmpcfg[0][7:0] {
		wildcard bins cfg_l000 = {8'b10011000};
		wildcard bins cfg_l001 = {8'b10011001};
		wildcard bins cfg_l011 = {8'b10011011};
		wildcard bins cfg_l100 = {8'b10011100};
		wildcard bins cfg_l101 = {8'b10011101};
		wildcard bins cfg_l111 = {8'b10011111};
	}

//-------------------------------------------------------

pmpcfgA_OFF: coverpoint {pmpcfg_a,pmp_hit} {
		wildcard bins OFF0  = {30'b????????????????????????????00_000000000000001};
		wildcard bins OFF1  = {30'b??????????????????????????00??_000000000000010};
		wildcard bins OFF2  = {30'b????????????????????????00????_000000000000100};
		wildcard bins OFF3  = {30'b??????????????????????00??????_000000000001000};
		wildcard bins OFF4  = {30'b????????????????????00????????_000000000010000};
		wildcard bins OFF5  = {30'b??????????????????00??????????_000000000100000};
		wildcard bins OFF6  = {30'b????????????????00????????????_000000001000000};
		wildcard bins OFF7  = {30'b??????????????00??????????????_000000010000000};
		wildcard bins OFF8  = {30'b????????????00????????????????_000000100000000};
		wildcard bins OFF9  = {30'b??????????00??????????????????_000001000000000};
		wildcard bins OFF10 = {30'b????????00????????????????????_000010000000000};
		wildcard bins OFF11 = {30'b??????00??????????????????????_000100000000000};
		wildcard bins OFF12 = {30'b????00????????????????????????_001000000000000};
		wildcard bins OFF13 = {30'b??00??????????????????????????_010000000000000};
		wildcard bins OFF14 = {30'b00????????????????????????????_100000000000000};
	}
	pmpcfgA_TOR: coverpoint {pmpcfg_a,pmp_hit} {
		wildcard bins TOR0  = {30'b????????????????????????????01_000000000000001};
		wildcard bins TOR1  = {30'b??????????????????????????01??_000000000000010};
		wildcard bins TOR2  = {30'b????????????????????????01????_000000000000100};
		wildcard bins TOR3  = {30'b??????????????????????01??????_000000000001000};
		wildcard bins TOR4  = {30'b????????????????????01????????_000000000010000};
		wildcard bins TOR5  = {30'b??????????????????01??????????_000000000100000};
		wildcard bins TOR6  = {30'b????????????????01????????????_000000001000000};
		wildcard bins TOR7  = {30'b??????????????01??????????????_000000010000000};
		wildcard bins TOR8  = {30'b????????????01????????????????_000000100000000};
		wildcard bins TOR9  = {30'b??????????01??????????????????_000001000000000};
		wildcard bins TOR10 = {30'b????????01????????????????????_000010000000000};
		wildcard bins TOR11 = {30'b??????01??????????????????????_000100000000000};
		wildcard bins TOR12 = {30'b????01????????????????????????_001000000000000};
		wildcard bins TOR13 = {30'b??01??????????????????????????_010000000000000};
		wildcard bins TOR14 = {30'b01????????????????????????????_100000000000000};
	}
	pmpcfgA_NA4: coverpoint {pmpcfg_a,pmp_hit} iff(`G==0){ //only fire these bins when G = 0
		wildcard bins NA40  = {30'b????????????????????????????10_000000000000001};
		wildcard bins NA41  = {30'b??????????????????????????10??_000000000000010};
		wildcard bins NA42  = {30'b????????????????????????10????_000000000000100};
		wildcard bins NA43  = {30'b??????????????????????10??????_000000000001000};
		wildcard bins NA44  = {30'b????????????????????10????????_000000000010000};
		wildcard bins NA45  = {30'b??????????????????10??????????_000000000100000};
		wildcard bins NA46  = {30'b????????????????10????????????_000000001000000};
		wildcard bins NA47  = {30'b??????????????10??????????????_000000010000000};
		wildcard bins NA48  = {30'b????????????10????????????????_000000100000000};
		wildcard bins NA49  = {30'b??????????10??????????????????_000001000000000};
		wildcard bins NA410 = {30'b????????10????????????????????_000010000000000};
		wildcard bins NA411 = {30'b??????10??????????????????????_000100000000000};
		wildcard bins NA412 = {30'b????10????????????????????????_001000000000000};
		wildcard bins NA413 = {30'b??10??????????????????????????_010000000000000};
		wildcard bins NA414 = {30'b10????????????????????????????_100000000000000};
	}
	pmpcfgA_NAPOT: coverpoint {pmpcfg_a,pmp_hit} {
		wildcard bins NAPOT0  = {30'b????????????????????????????11_000000000000001};
		wildcard bins NAPOT1  = {30'b??????????????????????????11??_000000000000010};
		wildcard bins NAPOT2  = {30'b????????????????????????11????_000000000000100};
		wildcard bins NAPOT3  = {30'b??????????????????????11??????_000000000001000};
		wildcard bins NAPOT4  = {30'b????????????????????11????????_000000000010000};
		wildcard bins NAPOT5  = {30'b??????????????????11??????????_000000000100000};
		wildcard bins NAPOT6  = {30'b????????????????11????????????_000000001000000};
		wildcard bins NAPOT7  = {30'b??????????????11??????????????_000000010000000};
		wildcard bins NAPOT8  = {30'b????????????11????????????????_000000100000000};
		wildcard bins NAPOT9  = {30'b??????????11??????????????????_000001000000000};
		wildcard bins NAPOT10 = {30'b????????11????????????????????_000010000000000};
		wildcard bins NAPOT11 = {30'b??????11??????????????????????_000100000000000};
		wildcard bins NAPOT12 = {30'b????11????????????????????????_001000000000000};
		wildcard bins NAPOT13 = {30'b??11??????????????????????????_010000000000000};
		wildcard bins NAPOT14 = {30'b11????????????????????????????_100000000000000};
	}

//-------------------------------------------------------

	RWXL000: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 0
		wildcard bins pmp0cfg_rwx000  = {75'b????????????????????????????00_??????????????0_??????????????0_000000000000001};
		wildcard bins pmp1cfg_rwx000  = {75'b??????????????????????????00??_?????????????0?_?????????????0?_000000000000010};
		wildcard bins pmp2cfg_rwx000  = {75'b????????????????????????00????_????????????0??_????????????0??_000000000000100};
		wildcard bins pmp3cfg_rwx000  = {75'b??????????????????????00??????_???????????0???_???????????0???_000000000001000};
		wildcard bins pmp4cfg_rwx000  = {75'b????????????????????00????????_??????????0????_??????????0????_000000000010000};
		wildcard bins pmp5cfg_rwx000  = {75'b??????????????????00??????????_?????????0?????_?????????0?????_000000000100000};
		wildcard bins pmp6cfg_rwx000  = {75'b????????????????00????????????_????????0??????_????????0??????_000000001000000};
		wildcard bins pmp7cfg_rwx000  = {75'b??????????????00??????????????_???????0???????_???????0???????_000000010000000};
		wildcard bins pmp8cfg_rwx000  = {75'b????????????00????????????????_??????0????????_??????0????????_000000100000000};
		wildcard bins pmp9cfg_rwx000  = {75'b??????????00??????????????????_?????0?????????_?????0?????????_000001000000000};
		wildcard bins pmp10cfg_rwx000 = {75'b????????00????????????????????_????0??????????_????0??????????_000010000000000};
		wildcard bins pmp11cfg_rwx000 = {75'b??????00??????????????????????_???0???????????_???0???????????_000100000000000};
		wildcard bins pmp12cfg_rwx000 = {75'b????00????????????????????????_??0????????????_??0????????????_001000000000000};
		wildcard bins pmp13cfg_rwx000 = {75'b??00??????????????????????????_?0?????????????_?0?????????????_010000000000000};
		wildcard bins pmp14cfg_rwx000 = {75'b00????????????????????????????_0??????????????_0??????????????_100000000000000};
	}

//-------------------------------------------------------

  legal_RWX_L_NAPOT: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = legal combinations, pmpcfg.L = 1 and pmpcfg.A = 3 for region pmp0
		wildcard bins pmp0cfg_rwx000  = {105'b????????????????????????????00_??????????????0_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp0cfg_rwx001  = {105'b????????????????????????????00_??????????????1_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp0cfg_rwx101  = {105'b????????????????????????????00_??????????????1_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp0cfg_rwx011  = {105'b????????????????????????????01_??????????????1_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp0cfg_rwx100  = {105'b????????????????????????????10_??????????????0_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp0cfg_rwx111  = {105'b????????????????????????????11_??????????????1_??????????????1_????????????????????????????11_000000000000001};
	}

//-------------------------------------------------------
  legal_RWX_L_NA4: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} iff(`G==0){ // pmpcfg.RWX = legal combinations, pmpcfg.L = 1 and pmpcfg.A = 2'b10 for region pmp0
		wildcard bins pmp0cfg_rwx000  = {105'b????????????????????????????00_??????????????0_??????????????1_????????????????????????????10_000000000000001};
		wildcard bins pmp0cfg_rwx001  = {105'b????????????????????????????00_??????????????1_??????????????1_????????????????????????????10_000000000000001};
		wildcard bins pmp0cfg_rwx101  = {105'b????????????????????????????00_??????????????1_??????????????1_????????????????????????????10_000000000000001};
		wildcard bins pmp0cfg_rwx011  = {105'b????????????????????????????01_??????????????1_??????????????1_????????????????????????????10_000000000000001};
		wildcard bins pmp0cfg_rwx100  = {105'b????????????????????????????10_??????????????0_??????????????1_????????????????????????????10_000000000000001};
		wildcard bins pmp0cfg_rwx111  = {105'b????????????????????????????11_??????????????1_??????????????1_????????????????????????????10_000000000000001};
	}

//-------------------------------------------------------
	RWXL001: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 1
		wildcard bins pmp0cfg_rwx000  = {75'b????????????????????????????00_??????????????0_??????????????1_000000000000001};
		wildcard bins pmp1cfg_rwx000  = {75'b??????????????????????????00??_?????????????0?_?????????????1?_000000000000010};
		wildcard bins pmp2cfg_rwx000  = {75'b????????????????????????00????_????????????0??_????????????1??_000000000000100};
		wildcard bins pmp3cfg_rwx000  = {75'b??????????????????????00??????_???????????0???_???????????1???_000000000001000};
		wildcard bins pmp4cfg_rwx000  = {75'b????????????????????00????????_??????????0????_??????????1????_000000000010000};
		wildcard bins pmp5cfg_rwx000  = {75'b??????????????????00??????????_?????????0?????_?????????1?????_000000000100000};
		wildcard bins pmp6cfg_rwx000  = {75'b????????????????00????????????_????????0??????_????????1??????_000000001000000};
		wildcard bins pmp7cfg_rwx000  = {75'b??????????????00??????????????_???????0???????_???????1???????_000000010000000};
		wildcard bins pmp8cfg_rwx000  = {75'b????????????00????????????????_??????0????????_??????1????????_000000100000000};
		wildcard bins pmp9cfg_rwx000  = {75'b??????????00??????????????????_?????0?????????_?????1?????????_000001000000000};
		wildcard bins pmp10cfg_rwx000 = {75'b????????00????????????????????_????0??????????_????1??????????_000010000000000};
		wildcard bins pmp11cfg_rwx000 = {75'b??????00??????????????????????_???0???????????_???1???????????_000100000000000};
		wildcard bins pmp12cfg_rwx000 = {75'b????00????????????????????????_??0????????????_??1????????????_001000000000000};
		wildcard bins pmp13cfg_rwx000 = {75'b??00??????????????????????????_?0?????????????_?1?????????????_010000000000000};
		wildcard bins pmp14cfg_rwx000 = {75'b00????????????????????????????_0??????????????_1??????????????_100000000000000};
	}

//-------------------------------------------------------

	X0: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x0   = {75'b??????????????0_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_x0   = {75'b?????????????0?_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_x0   = {75'b????????????0??_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_x0   = {75'b???????????0???_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_x0   = {75'b??????????0????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_x0   = {75'b?????????0?????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_x0   = {75'b????????0??????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_x0   = {75'b???????0???????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_x0   = {75'b??????0????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_x0   = {75'b?????0?????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_x0  = {75'b????0??????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_x0  = {75'b???0???????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_x0  = {75'b??0????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_x0  = {75'b?0?????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_x0  = {75'b0??????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	X1: coverpoint {pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.X = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_x1   = {75'b??????????????1_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_x1   = {75'b?????????????1?_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_x1   = {75'b????????????1??_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_x1   = {75'b???????????1???_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_x1   = {75'b??????????1????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_x1   = {75'b?????????1?????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_x1   = {75'b????????1??????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_x1   = {75'b???????1???????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_x1   = {75'b??????1????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_x1   = {75'b?????1?????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_x1  = {75'b????1??????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_x1  = {75'b???1???????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_x1  = {75'b??1????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_x1  = {75'b?1?????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_x1  = {75'b1??????????????_1??????????????_11????????????????????????????_100000000000000};
	}

//-------------------------------------------------------

	RW00: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 0, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw00   = {90'b????????????????????????????00_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw00   = {90'b??????????????????????????00??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw00   = {90'b????????????????????????00????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw00   = {90'b??????????????????????00??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw00   = {90'b????????????????????00????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw00   = {90'b??????????????????00??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw00   = {90'b????????????????00????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw00   = {90'b??????????????00??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw00   = {90'b????????????00????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw00   = {90'b??????????00??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw00  = {90'b????????00????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw00  = {90'b??????00??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw00  = {90'b????00????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw00  = {90'b??00??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw00  = {90'b00????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	RW11: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 3, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????11_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????11??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????11????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????11??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????11????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????11??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????11????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????11??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw11     = {90'b????????????11????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw11     = {90'b??????????11??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw11    = {90'b????????11????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw11    = {90'b??????11??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw11    = {90'b????11????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw11    = {90'b??11??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw11    = {90'b11????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

	RW10: coverpoint {pmpcfg_rw, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RW = 1, pmpcfg.L = 1 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rw11     = {90'b????????????????????????????01_??????????????1_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rw11     = {90'b??????????????????????????01??_?????????????1?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rw11     = {90'b????????????????????????01????_????????????1??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rw11     = {90'b??????????????????????01??????_???????????1???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rw11     = {90'b????????????????????01????????_??????????1????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rw11     = {90'b??????????????????01??????????_?????????1?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rw11     = {90'b????????????????01????????????_????????1??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rw11     = {90'b??????????????01??????????????_???????1???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rw11     = {90'b????????????01????????????????_??????1????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rw11     = {90'b??????????01??????????????????_?????1?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rw11    = {90'b????????01????????????????????_????1??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rw11    = {90'b??????01??????????????????????_???1???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rw11    = {90'b????01????????????????????????_??1????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rw11    = {90'b??01??????????????????????????_?1?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rw11    = {90'b01????????????????????????????_1??????????????_11????????????????????????????_100000000000000};
	}

//-------------------------------------------------------

	RWX000: coverpoint {pmpcfg_rw, pmpcfg_x, pmpcfg_l, pmpcfg_a, pmp_hit} { // pmpcfg.RWX = 0, pmpcfg.L = 0 and pmpcfg.A = 3
		wildcard bins pmp0cfg_rwx000  = {105'b????????????????????????????00_??????????????0_??????????????0_????????????????????????????11_000000000000001};
		wildcard bins pmp1cfg_rwx000  = {105'b??????????????????????????00??_?????????????0?_?????????????0?_??????????????????????????11??_000000000000010};
		wildcard bins pmp2cfg_rwx000  = {105'b????????????????????????00????_????????????0??_????????????0??_????????????????????????11????_000000000000100};
		wildcard bins pmp3cfg_rwx000  = {105'b??????????????????????00??????_???????????0???_???????????0???_??????????????????????11??????_000000000001000};
		wildcard bins pmp4cfg_rwx000  = {105'b????????????????????00????????_??????????0????_??????????0????_????????????????????11????????_000000000010000};
		wildcard bins pmp5cfg_rwx000  = {105'b??????????????????00??????????_?????????0?????_?????????0?????_??????????????????11??????????_000000000100000};
		wildcard bins pmp6cfg_rwx000  = {105'b????????????????00????????????_????????0??????_????????0??????_????????????????11????????????_000000001000000};
		wildcard bins pmp7cfg_rwx000  = {105'b??????????????00??????????????_???????0???????_???????0???????_??????????????11??????????????_000000010000000};
		wildcard bins pmp8cfg_rwx000  = {105'b????????????00????????????????_??????0????????_??????0????????_????????????11????????????????_000000100000000};
		wildcard bins pmp9cfg_rwx000  = {105'b??????????00??????????????????_?????0?????????_?????0?????????_??????????11??????????????????_000001000000000};
		wildcard bins pmp10cfg_rwx000 = {105'b????????00????????????????????_????0??????????_????0??????????_????????11????????????????????_000010000000000};
		wildcard bins pmp11cfg_rwx000 = {105'b??????00??????????????????????_???0???????????_???0???????????_??????11??????????????????????_000100000000000};
		wildcard bins pmp12cfg_rwx000 = {105'b????00????????????????????????_??0????????????_??0????????????_????11????????????????????????_001000000000000};
		wildcard bins pmp13cfg_rwx000 = {105'b??00??????????????????????????_?0?????????????_?0?????????????_??11??????????????????????????_010000000000000};
		wildcard bins pmp14cfg_rwx000 = {105'b00????????????????????????????_0??????????????_0??????????????_11????????????????????????????_100000000000000};
	}

//-------------------------------------------------------

	// Lock pmp_region_1 and check the writes on pmp_region_1 and pmp_region_0
	lock_checking: coverpoint pmpcfg_l[1] {
		bins region_locked = {1'b1};
		bins region_unlocked = {1'b0};
	}

	// Setting pmp_region_1 so incase of TOR we can check lock for pmp_region_0
	pmp_region: coverpoint pmpcfg[1][12:11] {
		bins OFF   = {2'b00};
		bins TOR   = {2'b01};
		bins NAPOT = {2'b11};
	}

	pmpcfg_xwr: coverpoint ins.prev.csr[12'h3A1][6:0] { // Region 1
		bins NAPOT_XWR = {7'b0011111};
	}

	lower_pmpcfg_xwr: coverpoint ins.prev.csr[12'h3A0][6:0] { // Region 0
		bins NAPOT_XWR = {7'b0000000};
	}

	pmpaddr: coverpoint ins.prev.csr[12'h3B1] { // Region 1
		bins hex_0x100 = {256};
	}

	rs1_val_for_pmpcfg: coverpoint ins.prev.rs1_val { // It will try to change pmpcfg_i-1 to 00000111
		bins pmpcfg_val = {7};
	}

	rs1_val_for_pmpaddr: coverpoint ins.prev.rs1_val { // It will try to change pmpaddr_i-1 to 0111 1111
		bins pmpaddr_val = {127};
	}

	write_pmp_csr: coverpoint ins.prev.insn {
		wildcard bins write_pmpaddr  = {32'b001110110001_00000_010_?????_1110011}; // Try to write value of x0 in pmpaddr[1]
		wildcard bins write_pmpcfg   = {32'b001110100001_00000_010_?????_1110011}; // Try to write value of x0 in pmpcfg[1]
	}

	write_lower_pmpaddr: coverpoint ins.prev.insn {
		wildcard bins write_pmpaddr  = {32'b001110110000_?????_010_?????_1110011}; // Try to write pmpaddr[0]
	}

	write_lower_pmpcfg: coverpoint ins.prev.insn {
		wildcard bins write_pmpcfg   = {32'b001110100000_?????_010_?????_1110011}; // Try to write pmpcfg[0]
	}

//-------------------------------------------------------

	cp_walk_rs1_pmpaddr: coverpoint ins.current.rs1_val {
		bins all_zeros = {0};
		bins all_ones = {-1};
		`ifdef XLEN32
			wildcard bins walking_ones_0  = {32'b00000000000000000000000000000001};
			wildcard bins walking_ones_1  = {32'b00000000000000000000000000000010};
			wildcard bins walking_ones_2  = {32'b00000000000000000000000000000100};
			wildcard bins walking_ones_3  = {32'b00000000000000000000000000001000};
			wildcard bins walking_ones_4  = {32'b00000000000000000000000000010000};
			wildcard bins walking_ones_5  = {32'b00000000000000000000000000100000};
			wildcard bins walking_ones_6  = {32'b00000000000000000000000001000000};
			wildcard bins walking_ones_7  = {32'b00000000000000000000000010000000};
			wildcard bins walking_ones_8  = {32'b00000000000000000000000100000000};
			wildcard bins walking_ones_9  = {32'b00000000000000000000001000000000};
			wildcard bins walking_ones_10 = {32'b00000000000000000000010000000000};
			wildcard bins walking_ones_11 = {32'b00000000000000000000100000000000};
			wildcard bins walking_ones_12 = {32'b00000000000000000001000000000000};
			wildcard bins walking_ones_13 = {32'b00000000000000000010000000000000};
			wildcard bins walking_ones_14 = {32'b00000000000000000100000000000000};
			wildcard bins walking_ones_15 = {32'b00000000000000001000000000000000};
			wildcard bins walking_ones_16 = {32'b00000000000000010000000000000000};
			wildcard bins walking_ones_17 = {32'b00000000000000100000000000000000};
			wildcard bins walking_ones_18 = {32'b00000000000001000000000000000000};
			wildcard bins walking_ones_19 = {32'b00000000000010000000000000000000};
			wildcard bins walking_ones_20 = {32'b00000000000100000000000000000000};
			wildcard bins walking_ones_21 = {32'b00000000001000000000000000000000};
			wildcard bins walking_ones_22 = {32'b00000000010000000000000000000000};
			wildcard bins walking_ones_23 = {32'b00000000100000000000000000000000};
			wildcard bins walking_ones_24 = {32'b00000001000000000000000000000000};
			wildcard bins walking_ones_25 = {32'b00000010000000000000000000000000};
			wildcard bins walking_ones_26 = {32'b00000100000000000000000000000000};
			wildcard bins walking_ones_27 = {32'b00001000000000000000000000000000};
			wildcard bins walking_ones_28 = {32'b00010000000000000000000000000000};
			wildcard bins walking_ones_29 = {32'b00100000000000000000000000000000};
			wildcard bins walking_ones_30 = {32'b01000000000000000000000000000000};
			wildcard bins walking_ones_31 = {32'b10000000000000000000000000000000};
		`endif
		`ifdef XLEN64
			wildcard bins walking_ones_0  = {64'b??????????000000000000000000000000000000000000000000000000000001};
			wildcard bins walking_ones_1  = {64'b??????????000000000000000000000000000000000000000000000000000010};
			wildcard bins walking_ones_2  = {64'b??????????000000000000000000000000000000000000000000000000000100};
			wildcard bins walking_ones_3  = {64'b??????????000000000000000000000000000000000000000000000000001000};
			wildcard bins walking_ones_4  = {64'b??????????000000000000000000000000000000000000000000000000010000};
			wildcard bins walking_ones_5  = {64'b??????????000000000000000000000000000000000000000000000000100000};
			wildcard bins walking_ones_6  = {64'b??????????000000000000000000000000000000000000000000000001000000};
			wildcard bins walking_ones_7  = {64'b??????????000000000000000000000000000000000000000000000010000000};
			wildcard bins walking_ones_8  = {64'b??????????000000000000000000000000000000000000000000000100000000};
			wildcard bins walking_ones_9  = {64'b??????????000000000000000000000000000000000000000000001000000000};
			wildcard bins walking_ones_10 = {64'b??????????000000000000000000000000000000000000000000010000000000};
			wildcard bins walking_ones_11 = {64'b??????????000000000000000000000000000000000000000000100000000000};
			wildcard bins walking_ones_12 = {64'b??????????000000000000000000000000000000000000000001000000000000};
			wildcard bins walking_ones_13 = {64'b??????????000000000000000000000000000000000000000010000000000000};
			wildcard bins walking_ones_14 = {64'b??????????000000000000000000000000000000000000000100000000000000};
			wildcard bins walking_ones_15 = {64'b??????????000000000000000000000000000000000000001000000000000000};
			wildcard bins walking_ones_16 = {64'b??????????000000000000000000000000000000000000010000000000000000};
			wildcard bins walking_ones_17 = {64'b??????????000000000000000000000000000000000000100000000000000000};
			wildcard bins walking_ones_18 = {64'b??????????000000000000000000000000000000000001000000000000000000};
			wildcard bins walking_ones_19 = {64'b??????????000000000000000000000000000000000010000000000000000000};
			wildcard bins walking_ones_20 = {64'b??????????000000000000000000000000000000000100000000000000000000};
			wildcard bins walking_ones_21 = {64'b??????????000000000000000000000000000000001000000000000000000000};
			wildcard bins walking_ones_22 = {64'b??????????000000000000000000000000000000010000000000000000000000};
			wildcard bins walking_ones_23 = {64'b??????????000000000000000000000000000000100000000000000000000000};
			wildcard bins walking_ones_24 = {64'b??????????000000000000000000000000000001000000000000000000000000};
			wildcard bins walking_ones_25 = {64'b??????????000000000000000000000000000010000000000000000000000000};
			wildcard bins walking_ones_26 = {64'b??????????000000000000000000000000000100000000000000000000000000};
			wildcard bins walking_ones_27 = {64'b??????????000000000000000000000000001000000000000000000000000000};
			wildcard bins walking_ones_28 = {64'b??????????000000000000000000000000010000000000000000000000000000};
			wildcard bins walking_ones_29 = {64'b??????????000000000000000000000000100000000000000000000000000000};
			wildcard bins walking_ones_30 = {64'b??????????000000000000000000000001000000000000000000000000000000};
			wildcard bins walking_ones_31 = {64'b??????????000000000000000000000010000000000000000000000000000000};
			wildcard bins walking_ones_32 = {64'b??????????000000000000000000000100000000000000000000000000000000};
			wildcard bins walking_ones_33 = {64'b??????????000000000000000000001000000000000000000000000000000000};
			wildcard bins walking_ones_34 = {64'b??????????000000000000000000010000000000000000000000000000000000};
			wildcard bins walking_ones_35 = {64'b??????????000000000000000000100000000000000000000000000000000000};
			wildcard bins walking_ones_36 = {64'b??????????000000000000000001000000000000000000000000000000000000};
			wildcard bins walking_ones_37 = {64'b??????????000000000000000010000000000000000000000000000000000000};
			wildcard bins walking_ones_38 = {64'b??????????000000000000000100000000000000000000000000000000000000};
			wildcard bins walking_ones_39 = {64'b??????????000000000000001000000000000000000000000000000000000000};
			wildcard bins walking_ones_40 = {64'b??????????000000000000010000000000000000000000000000000000000000};
			wildcard bins walking_ones_41 = {64'b??????????000000000000100000000000000000000000000000000000000000};
			wildcard bins walking_ones_42 = {64'b??????????000000000001000000000000000000000000000000000000000000};
			wildcard bins walking_ones_43 = {64'b??????????000000000010000000000000000000000000000000000000000000};
			wildcard bins walking_ones_44 = {64'b??????????000000000100000000000000000000000000000000000000000000};
			wildcard bins walking_ones_45 = {64'b??????????000000001000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_46 = {64'b??????????000000010000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_47 = {64'b??????????000000100000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_48 = {64'b??????????000001000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_49 = {64'b??????????000010000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_50 = {64'b??????????000100000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_51 = {64'b??????????001000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_52 = {64'b??????????010000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_53 = {64'b??????????100000000000000000000000000000000000000000000000000000};
		`endif
	}

	cp_walk_rs1_pmpcfg: coverpoint ins.current.rs1_val {
		`ifdef XLEN32
			wildcard bins walking_ones_0  = {32'b00000000000000000000000000000001};
			wildcard bins walking_ones_1  = {32'b00000000000000000000000000000010};
			wildcard bins walking_ones_2  = {32'b00000000000000000000000000000100};
			wildcard bins walking_ones_3  = {32'b00000000000000000000000000001000};
			wildcard bins walking_ones_4  = {32'b00000000000000000000000000010000};
			wildcard bins walking_ones_5  = {32'b00000000000000000000000000100000};
			wildcard bins walking_ones_6  = {32'b00000000000000000000000001000000};
			wildcard bins walking_ones_7  = {32'b00000000000000000000000010000000};
			wildcard bins walking_ones_8  = {32'b00000000000000000000000100000000};
			wildcard bins walking_ones_9  = {32'b00000000000000000000001000000000};
			wildcard bins walking_ones_10 = {32'b00000000000000000000010000000000};
			wildcard bins walking_ones_11 = {32'b00000000000000000000100000000000};
			wildcard bins walking_ones_12 = {32'b00000000000000000001000000000000};
			wildcard bins walking_ones_13 = {32'b00000000000000000010000000000000};
			wildcard bins walking_ones_14 = {32'b00000000000000000100000000000000};
			wildcard bins walking_ones_15 = {32'b00000000000000001000000000000000};
			wildcard bins walking_ones_16 = {32'b00000000000000010000000000000000};
			wildcard bins walking_ones_17 = {32'b00000000000000100000000000000000};
			wildcard bins walking_ones_18 = {32'b00000000000001000000000000000000};
			wildcard bins walking_ones_19 = {32'b00000000000010000000000000000000};
			wildcard bins walking_ones_20 = {32'b00000000000100000000000000000000};
			wildcard bins walking_ones_21 = {32'b00000000001000000000000000000000};
			wildcard bins walking_ones_22 = {32'b00000000010000000000000000000000};
			wildcard bins walking_ones_23 = {32'b00000000100000000000000000000000};
			wildcard bins walking_ones_24 = {32'b00000001000000000000000000000000};
			wildcard bins walking_ones_25 = {32'b00000010000000000000000000000000};
			wildcard bins walking_ones_26 = {32'b00000100000000000000000000000000};
			wildcard bins walking_ones_27 = {32'b00001000000000000000000000000000};
			wildcard bins walking_ones_28 = {32'b00010000000000000000000000000000};
			wildcard bins walking_ones_29 = {32'b00100000000000000000000000000000};
			wildcard bins walking_ones_30 = {32'b01000000000000000000000000000000};
			wildcard bins walking_ones_31 = {32'b10000000000000000000000000000000};
		`endif
		`ifdef XLEN64
			wildcard bins walking_ones_0  = {64'b0000000000000000000000000000000000000000000000000000000000000001};
			wildcard bins walking_ones_1  = {64'b0000000000000000000000000000000000000000000000000000000000000010};
			wildcard bins walking_ones_2  = {64'b0000000000000000000000000000000000000000000000000000000000000100};
			wildcard bins walking_ones_3  = {64'b0000000000000000000000000000000000000000000000000000000000001000};
			wildcard bins walking_ones_4  = {64'b0000000000000000000000000000000000000000000000000000000000010000};
			wildcard bins walking_ones_5  = {64'b0000000000000000000000000000000000000000000000000000000000100000};
			wildcard bins walking_ones_6  = {64'b0000000000000000000000000000000000000000000000000000000001000000};
			wildcard bins walking_ones_7  = {64'b0000000000000000000000000000000000000000000000000000000010000000};
			wildcard bins walking_ones_8  = {64'b0000000000000000000000000000000000000000000000000000000100000000};
			wildcard bins walking_ones_9  = {64'b0000000000000000000000000000000000000000000000000000001000000000};
			wildcard bins walking_ones_10 = {64'b0000000000000000000000000000000000000000000000000000010000000000};
			wildcard bins walking_ones_11 = {64'b0000000000000000000000000000000000000000000000000000100000000000};
			wildcard bins walking_ones_12 = {64'b0000000000000000000000000000000000000000000000000001000000000000};
			wildcard bins walking_ones_13 = {64'b0000000000000000000000000000000000000000000000000010000000000000};
			wildcard bins walking_ones_14 = {64'b0000000000000000000000000000000000000000000000000100000000000000};
			wildcard bins walking_ones_15 = {64'b0000000000000000000000000000000000000000000000001000000000000000};
			wildcard bins walking_ones_16 = {64'b0000000000000000000000000000000000000000000000010000000000000000};
			wildcard bins walking_ones_17 = {64'b0000000000000000000000000000000000000000000000100000000000000000};
			wildcard bins walking_ones_18 = {64'b0000000000000000000000000000000000000000000001000000000000000000};
			wildcard bins walking_ones_19 = {64'b0000000000000000000000000000000000000000000010000000000000000000};
			wildcard bins walking_ones_20 = {64'b0000000000000000000000000000000000000000000100000000000000000000};
			wildcard bins walking_ones_21 = {64'b0000000000000000000000000000000000000000001000000000000000000000};
			wildcard bins walking_ones_22 = {64'b0000000000000000000000000000000000000000010000000000000000000000};
			wildcard bins walking_ones_23 = {64'b0000000000000000000000000000000000000000100000000000000000000000};
			wildcard bins walking_ones_24 = {64'b0000000000000000000000000000000000000001000000000000000000000000};
			wildcard bins walking_ones_25 = {64'b0000000000000000000000000000000000000010000000000000000000000000};
			wildcard bins walking_ones_26 = {64'b0000000000000000000000000000000000000100000000000000000000000000};
			wildcard bins walking_ones_27 = {64'b0000000000000000000000000000000000001000000000000000000000000000};
			wildcard bins walking_ones_28 = {64'b0000000000000000000000000000000000010000000000000000000000000000};
			wildcard bins walking_ones_29 = {64'b0000000000000000000000000000000000100000000000000000000000000000};
			wildcard bins walking_ones_30 = {64'b0000000000000000000000000000000001000000000000000000000000000000};
			wildcard bins walking_ones_31 = {64'b0000000000000000000000000000000010000000000000000000000000000000};
			wildcard bins walking_ones_32 = {64'b0000000000000000000000000000000100000000000000000000000000000000};
			wildcard bins walking_ones_33 = {64'b0000000000000000000000000000001000000000000000000000000000000000};
			wildcard bins walking_ones_34 = {64'b0000000000000000000000000000010000000000000000000000000000000000};
			wildcard bins walking_ones_35 = {64'b0000000000000000000000000000100000000000000000000000000000000000};
			wildcard bins walking_ones_36 = {64'b0000000000000000000000000001000000000000000000000000000000000000};
			wildcard bins walking_ones_37 = {64'b0000000000000000000000000010000000000000000000000000000000000000};
			wildcard bins walking_ones_38 = {64'b0000000000000000000000000100000000000000000000000000000000000000};
			wildcard bins walking_ones_39 = {64'b0000000000000000000000001000000000000000000000000000000000000000};
			wildcard bins walking_ones_40 = {64'b0000000000000000000000010000000000000000000000000000000000000000};
			wildcard bins walking_ones_41 = {64'b0000000000000000000000100000000000000000000000000000000000000000};
			wildcard bins walking_ones_42 = {64'b0000000000000000000001000000000000000000000000000000000000000000};
			wildcard bins walking_ones_43 = {64'b0000000000000000000010000000000000000000000000000000000000000000};
			wildcard bins walking_ones_44 = {64'b0000000000000000000100000000000000000000000000000000000000000000};
			wildcard bins walking_ones_45 = {64'b0000000000000000001000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_46 = {64'b0000000000000000010000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_47 = {64'b0000000000000000100000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_48 = {64'b0000000000000001000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_49 = {64'b0000000000000010000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_50 = {64'b0000000000000100000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_51 = {64'b0000000000001000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_52 = {64'b0000000000010000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_53 = {64'b0000000000100000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_54 = {64'b0000000001000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_55 = {64'b0000000010000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_56 = {64'b0000000100000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_57 = {64'b0000001000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_58 = {64'b0000010000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_59 = {64'b0000100000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_60 = {64'b0001000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_61 = {64'b0010000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_62 = {64'b0100000000000000000000000000000000000000000000000000000000000000};
			wildcard bins walking_ones_63 = {64'b1000000000000000000000000000000000000000000000000000000000000000};
		`endif
	}

	cp_zero_rs1: coverpoint ins.current.rs1_val {
		bins rs1_val = {0};
	}

	csrrw: coverpoint ins.current.insn {
		wildcard bins write_pmp_csr  = {32'b????????????_?????_010_?????_1110011}; // Try to write pmpaddr or pmpcfg
	}

	legal_pmpaddr_entries: coverpoint ins.current.insn[31:20] {
		bins pmpaddr0   = {12'h3B0};
		bins pmpaddr1   = {12'h3B1};
		bins pmpaddr2   = {12'h3B2};
		bins pmpaddr3   = {12'h3B3};
		bins pmpaddr4   = {12'h3B4};
		bins pmpaddr5   = {12'h3B5};
		bins pmpaddr6   = {12'h3B6};
		bins pmpaddr7   = {12'h3B7};
		bins pmpaddr8   = {12'h3B8};
		bins pmpaddr9   = {12'h3B9};
		bins pmpaddr10  = {12'h3BA};
		bins pmpaddr11  = {12'h3BB};
		bins pmpaddr12  = {12'h3BC};
		bins pmpaddr13  = {12'h3BD};
		bins pmpaddr14  = {12'h3BE};
		bins pmpaddr15  = {12'h3BF};
		`ifdef PMP_64
			bins pmpaddr16  = {12'h3C0};
			bins pmpaddr17  = {12'h3C1};
			bins pmpaddr18  = {12'h3C2};
			bins pmpaddr19  = {12'h3C3};
			bins pmpaddr20  = {12'h3C4};
			bins pmpaddr21  = {12'h3C5};
			bins pmpaddr22  = {12'h3C6};
			bins pmpaddr23  = {12'h3C7};
			bins pmpaddr24  = {12'h3C8};
			bins pmpaddr25  = {12'h3C9};
			bins pmpaddr26  = {12'h3CA};
			bins pmpaddr27  = {12'h3CB};
			bins pmpaddr28  = {12'h3CC};
			bins pmpaddr29  = {12'h3CD};
			bins pmpaddr30  = {12'h3CE};
			bins pmpaddr31  = {12'h3CF};
			bins pmpaddr32  = {12'h3D0};
			bins pmpaddr33  = {12'h3D1};
			bins pmpaddr34  = {12'h3D2};
			bins pmpaddr35  = {12'h3D3};
			bins pmpaddr36  = {12'h3D4};
			bins pmpaddr37  = {12'h3D5};
			bins pmpaddr38  = {12'h3D6};
			bins pmpaddr39  = {12'h3D7};
			bins pmpaddr40  = {12'h3D8};
			bins pmpaddr41  = {12'h3D9};
			bins pmpaddr42  = {12'h3DA};
			bins pmpaddr43  = {12'h3DB};
			bins pmpaddr44  = {12'h3DC};
			bins pmpaddr45  = {12'h3DD};
			bins pmpaddr46  = {12'h3DE};
			bins pmpaddr47  = {12'h3DF};
			bins pmpaddr48  = {12'h3E0};
			bins pmpaddr49  = {12'h3E1};
			bins pmpaddr50  = {12'h3E2};
			bins pmpaddr51  = {12'h3E3};
			bins pmpaddr52  = {12'h3E4};
			bins pmpaddr53  = {12'h3E5};
			bins pmpaddr54  = {12'h3E6};
			bins pmpaddr55  = {12'h3E7};
			bins pmpaddr56  = {12'h3E8};
			bins pmpaddr57  = {12'h3E9};
			bins pmpaddr58  = {12'h3EA};
			bins pmpaddr59  = {12'h3EB};
			bins pmpaddr60  = {12'h3EC};
			bins pmpaddr61  = {12'h3ED};
			bins pmpaddr62  = {12'h3EE};
			bins pmpaddr63  = {12'h3EF};
		`endif
	}

	legal_pmpcfg_entries_even: coverpoint ins.current.insn[31:20] { 	// For writing walking ones in even PMPCFGs
		bins pmpcfg0   = {12'h3A0};
		bins pmpcfg2   = {12'h3A2};
		`ifdef PMP_64
			bins pmpcfg4   = {12'h3A4};
			bins pmpcfg6   = {12'h3A6};
			bins pmpcfg8   = {12'h3A8};
			bins pmpcfg10  = {12'h3AA};
			bins pmpcfg12  = {12'h3AC};
			bins pmpcfg14  = {12'h3AE};
		`endif
	}

	legal_pmpcfg_entries_odd: coverpoint ins.current.insn[31:20] { 	// For writing zero in odd PMPCFGs
		bins pmpcfg1   = {12'h3A1};
		bins pmpcfg3   = {12'h3A3};
		`ifdef PMP_64
			bins pmpcfg5   = {12'h3A5};
			bins pmpcfg7   = {12'h3A7};
			bins pmpcfg9   = {12'h3A9};
			bins pmpcfg11  = {12'h3AB};
			bins pmpcfg13  = {12'h3AD};
			bins pmpcfg15  = {12'h3AF};
		`endif
	}
//-------------------------------------------------------

	pmp64: coverpoint {pmpcfg_L, pmpcfg_X, pmpcfg_RW, pmp_HIT} {
		wildcard bins pmp15cfg = {240'b???????????????????????????????????????????????1_???????????????????????????????????????????????1_??????????????????????????????????????????????????????????????????????????????????????????????01_000000000000000000000000000000000000000000000001};
		wildcard bins pmp16cfg = {240'b??????????????????????????????????????????????1?_??????????????????????????????????????????????1?_????????????????????????????????????????????????????????????????????????????????????????????01??_000000000000000000000000000000000000000000000010};
		wildcard bins pmp17cfg = {240'b?????????????????????????????????????????????1??_?????????????????????????????????????????????1??_??????????????????????????????????????????????????????????????????????????????????????????01????_000000000000000000000000000000000000000000000100};
		wildcard bins pmp18cfg = {240'b????????????????????????????????????????????1???_????????????????????????????????????????????1???_????????????????????????????????????????????????????????????????????????????????????????01??????_000000000000000000000000000000000000000000001000};
		wildcard bins pmp19cfg = {240'b???????????????????????????????????????????1????_???????????????????????????????????????????1????_??????????????????????????????????????????????????????????????????????????????????????01????????_000000000000000000000000000000000000000000010000};
		wildcard bins pmp20cfg = {240'b??????????????????????????????????????????1?????_??????????????????????????????????????????1?????_????????????????????????????????????????????????????????????????????????????????????01??????????_000000000000000000000000000000000000000000100000};
		wildcard bins pmp21cfg = {240'b?????????????????????????????????????????1??????_?????????????????????????????????????????1??????_??????????????????????????????????????????????????????????????????????????????????01????????????_000000000000000000000000000000000000000001000000};
		wildcard bins pmp22cfg = {240'b????????????????????????????????????????1???????_????????????????????????????????????????1???????_????????????????????????????????????????????????????????????????????????????????01??????????????_000000000000000000000000000000000000000010000000};
		wildcard bins pmp23cfg = {240'b???????????????????????????????????????1????????_???????????????????????????????????????1????????_??????????????????????????????????????????????????????????????????????????????01????????????????_000000000000000000000000000000000000000100000000};
		wildcard bins pmp24cfg = {240'b??????????????????????????????????????1?????????_??????????????????????????????????????1?????????_????????????????????????????????????????????????????????????????????????????01??????????????????_000000000000000000000000000000000000001000000000};
		wildcard bins pmp25cfg = {240'b?????????????????????????????????????1??????????_?????????????????????????????????????1??????????_??????????????????????????????????????????????????????????????????????????01????????????????????_000000000000000000000000000000000000010000000000};
		wildcard bins pmp26cfg = {240'b????????????????????????????????????1???????????_????????????????????????????????????1???????????_????????????????????????????????????????????????????????????????????????01??????????????????????_000000000000000000000000000000000000100000000000};
		wildcard bins pmp27cfg = {240'b???????????????????????????????????1????????????_???????????????????????????????????1????????????_??????????????????????????????????????????????????????????????????????01????????????????????????_000000000000000000000000000000000001000000000000};
		wildcard bins pmp28cfg = {240'b??????????????????????????????????1?????????????_??????????????????????????????????1?????????????_????????????????????????????????????????????????????????????????????01??????????????????????????_000000000000000000000000000000000010000000000000};
		wildcard bins pmp29cfg = {240'b?????????????????????????????????1??????????????_?????????????????????????????????1??????????????_??????????????????????????????????????????????????????????????????01????????????????????????????_000000000000000000000000000000000100000000000000};
		wildcard bins pmp30cfg = {240'b????????????????????????????????1???????????????_????????????????????????????????1???????????????_????????????????????????????????????????????????????????????????01??????????????????????????????_000000000000000000000000000000001000000000000000};
		wildcard bins pmp31cfg = {240'b???????????????????????????????1????????????????_???????????????????????????????1????????????????_??????????????????????????????????????????????????????????????01????????????????????????????????_000000000000000000000000000000010000000000000000};
		wildcard bins pmp32cfg = {240'b??????????????????????????????1?????????????????_??????????????????????????????1?????????????????_????????????????????????????????????????????????????????????01??????????????????????????????????_000000000000000000000000000000100000000000000000};
		wildcard bins pmp33cfg = {240'b?????????????????????????????1??????????????????_?????????????????????????????1??????????????????_??????????????????????????????????????????????????????????01????????????????????????????????????_000000000000000000000000000001000000000000000000};
		wildcard bins pmp34cfg = {240'b????????????????????????????1???????????????????_????????????????????????????1???????????????????_????????????????????????????????????????????????????????01??????????????????????????????????????_000000000000000000000000000010000000000000000000};
		wildcard bins pmp35cfg = {240'b???????????????????????????1????????????????????_???????????????????????????1????????????????????_??????????????????????????????????????????????????????01????????????????????????????????????????_000000000000000000000000000100000000000000000000};
		wildcard bins pmp36cfg = {240'b??????????????????????????1?????????????????????_??????????????????????????1?????????????????????_????????????????????????????????????????????????????01??????????????????????????????????????????_000000000000000000000000001000000000000000000000};
		wildcard bins pmp37cfg = {240'b?????????????????????????1??????????????????????_?????????????????????????1??????????????????????_??????????????????????????????????????????????????01????????????????????????????????????????????_000000000000000000000000010000000000000000000000};
		wildcard bins pmp38cfg = {240'b????????????????????????1???????????????????????_????????????????????????1???????????????????????_????????????????????????????????????????????????01??????????????????????????????????????????????_000000000000000000000000100000000000000000000000};
		wildcard bins pmp39cfg = {240'b???????????????????????1????????????????????????_???????????????????????1????????????????????????_??????????????????????????????????????????????01????????????????????????????????????????????????_000000000000000000000001000000000000000000000000};
		wildcard bins pmp40cfg = {240'b??????????????????????1?????????????????????????_??????????????????????1?????????????????????????_????????????????????????????????????????????01??????????????????????????????????????????????????_000000000000000000000010000000000000000000000000};
		wildcard bins pmp41cfg = {240'b?????????????????????1??????????????????????????_?????????????????????1??????????????????????????_??????????????????????????????????????????01????????????????????????????????????????????????????_000000000000000000000100000000000000000000000000};
		wildcard bins pmp42cfg = {240'b????????????????????1???????????????????????????_????????????????????1???????????????????????????_????????????????????????????????????????01??????????????????????????????????????????????????????_000000000000000000001000000000000000000000000000};
		wildcard bins pmp43cfg = {240'b???????????????????1????????????????????????????_???????????????????1????????????????????????????_??????????????????????????????????????01????????????????????????????????????????????????????????_000000000000000000010000000000000000000000000000};
		wildcard bins pmp44cfg = {240'b??????????????????1?????????????????????????????_??????????????????1?????????????????????????????_????????????????????????????????????01??????????????????????????????????????????????????????????_000000000000000000100000000000000000000000000000};
		wildcard bins pmp45cfg = {240'b?????????????????1??????????????????????????????_?????????????????1??????????????????????????????_??????????????????????????????????01????????????????????????????????????????????????????????????_000000000000000001000000000000000000000000000000};
		wildcard bins pmp46cfg = {240'b????????????????1???????????????????????????????_????????????????1???????????????????????????????_????????????????????????????????01??????????????????????????????????????????????????????????????_000000000000000010000000000000000000000000000000};
		wildcard bins pmp47cfg = {240'b???????????????1????????????????????????????????_???????????????1????????????????????????????????_??????????????????????????????01????????????????????????????????????????????????????????????????_000000000000000100000000000000000000000000000000};
		wildcard bins pmp48cfg = {240'b??????????????1?????????????????????????????????_??????????????1?????????????????????????????????_????????????????????????????01??????????????????????????????????????????????????????????????????_000000000000001000000000000000000000000000000000};
		wildcard bins pmp49cfg = {240'b?????????????1??????????????????????????????????_?????????????1??????????????????????????????????_??????????????????????????01????????????????????????????????????????????????????????????????????_000000000000010000000000000000000000000000000000};
		wildcard bins pmp50cfg = {240'b????????????1???????????????????????????????????_????????????1???????????????????????????????????_????????????????????????01??????????????????????????????????????????????????????????????????????_000000000000100000000000000000000000000000000000};
		wildcard bins pmp51cfg = {240'b???????????1????????????????????????????????????_???????????1????????????????????????????????????_??????????????????????01????????????????????????????????????????????????????????????????????????_000000000001000000000000000000000000000000000000};
		wildcard bins pmp52cfg = {240'b??????????1?????????????????????????????????????_??????????1?????????????????????????????????????_????????????????????01??????????????????????????????????????????????????????????????????????????_000000000010000000000000000000000000000000000000};
		wildcard bins pmp53cfg = {240'b?????????1??????????????????????????????????????_?????????1??????????????????????????????????????_??????????????????01????????????????????????????????????????????????????????????????????????????_000000000100000000000000000000000000000000000000};
		wildcard bins pmp54cfg = {240'b????????1???????????????????????????????????????_????????1???????????????????????????????????????_????????????????01??????????????????????????????????????????????????????????????????????????????_000000001000000000000000000000000000000000000000};
		wildcard bins pmp55cfg = {240'b???????1????????????????????????????????????????_???????1????????????????????????????????????????_??????????????01????????????????????????????????????????????????????????????????????????????????_000000010000000000000000000000000000000000000000};
		wildcard bins pmp56cfg = {240'b??????1?????????????????????????????????????????_??????1?????????????????????????????????????????_????????????01??????????????????????????????????????????????????????????????????????????????????_000000100000000000000000000000000000000000000000};
		wildcard bins pmp57cfg = {240'b?????1??????????????????????????????????????????_?????1??????????????????????????????????????????_??????????01????????????????????????????????????????????????????????????????????????????????????_000001000000000000000000000000000000000000000000};
		wildcard bins pmp58cfg = {240'b????1???????????????????????????????????????????_????1???????????????????????????????????????????_????????01??????????????????????????????????????????????????????????????????????????????????????_000010000000000000000000000000000000000000000000};
		wildcard bins pmp59cfg = {240'b???1????????????????????????????????????????????_???1????????????????????????????????????????????_??????01????????????????????????????????????????????????????????????????????????????????????????_000100000000000000000000000000000000000000000000};
		wildcard bins pmp61cfg = {240'b??1?????????????????????????????????????????????_??1?????????????????????????????????????????????_????01??????????????????????????????????????????????????????????????????????????????????????????_001000000000000000000000000000000000000000000000};
		wildcard bins pmp62cfg = {240'b?1??????????????????????????????????????????????_?1??????????????????????????????????????????????_??01????????????????????????????????????????????????????????????????????????????????????????????_010000000000000000000000000000000000000000000000};
		wildcard bins pmp63cfg = {240'b1???????????????????????????????????????????????_1???????????????????????????????????????????????_01??????????????????????????????????????????????????????????????????????????????????????????????_100000000000000000000000000000000000000000000000};
	}

//-------------------------------------------------------

	cp_cfg_X: cross priv_mode_m, legal_lxwr, exec_instr, standard_region, addr_in_region ;
	cp_cfg_R: cross priv_mode_m, legal_lxwr, read_instr, standard_region, addr_in_region ;
	cp_cfg_W: cross priv_mode_m, legal_lxwr, write_instr, standard_region, addr_in_region ;

	cp_cfg_X1_all: cross priv_mode_m, exec_instr, X1, addr_in_region ;
	cp_cfg_X0_all: cross priv_mode_m, exec_instr, X0, addr_in_region ;

	cp_cfg_Rw00_all: cross priv_mode_m, read_instr, RW00, addr_in_region ;
	cp_cfg_Rw10_all: cross priv_mode_m, read_instr, RW10, addr_in_region ;
	cp_cfg_Rw11_all: cross priv_mode_m, read_instr, RW11, addr_in_region ;
	cp_cfg_rW00_all: cross priv_mode_m, write_instr, RW00, addr_in_region ;
	cp_cfg_rW10_all: cross priv_mode_m, write_instr, RW10, addr_in_region ;
	cp_cfg_rW11_all: cross priv_mode_m, write_instr, RW11, addr_in_region ;

	cp_cfg_L_access_exec: cross priv_mode_m, exec_instr, RWX000, addr_in_region ;
	cp_cfg_L_access_read: cross priv_mode_m, read_instr, RWX000, addr_in_region ;
	cp_cfg_L_access_write: cross priv_mode_m, write_instr, RWX000, addr_in_region ;

	cp_cfg_L_modify: cross priv_mode_m, lock_checking, pmp_region, write_pmp_csr, pmpcfg_xwr, pmpaddr ;
	// If pmpcfg.A = TOR and pmpcfg.L = 1, pmpaddr_i-1 will be unchange but not pmpcfg_i-1.

  cp_cfg_L_modify_TOR_pmpaddr: cross priv_mode_m, lock_checking, pmp_region, write_lower_pmpaddr, rs1_val_for_pmpaddr, lower_pmpcfg_xwr, pmpaddr ;
	cp_cfg_L_modify_TOR_pmpcfg: cross priv_mode_m, lock_checking, pmp_region, write_lower_pmpcfg, rs1_val_for_pmpcfg, lower_pmpcfg_xwr, pmpaddr ;

	cp_pmpaddr_walk: cross priv_mode_m, cp_walk_rs1, csrrw, legal_pmpaddr_entries;
	cp_pmpcfg_walk: cross priv_mode_m, cp_walk_rs1, csrrw, legal_pmpcfg_entries;

	cp_cfg_A_OFF_allr : cross pmpcfgA_OFF, RWXL001, read_instr, addr_in_region;
	cp_cfg_A_OFF_allw : cross pmpcfgA_OFF, RWXL001, write_instr, addr_in_region;
	cp_cfg_A_OFF_allx : cross pmpcfgA_OFF, RWXL001, exec_instr, addr_in_region;

	cp_cfg_A_napot_all: cross pmpcfgA_NAPOT, RWXL001, read_instr_lw, addr_offset{
		ignore_bins ig5  = binsof(addr_offset.above_base);
		ignore_bins ig6  = binsof(addr_offset.highest_word);
	}

	cp_cfg_A_napot_x : cross legal_RWX_L_NAPOT, addr_offset, exec_instr{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}
	cp_cfg_A_napot_r : cross legal_RWX_L_NAPOT, addr_offset, read_instr_lw{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}
	cp_cfg_A_napot_w : cross legal_RWX_L_NAPOT, addr_offset, write_instr_sw{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}

	cp_cfg_A_na4_x : cross legal_RWX_L_NA4, addr_offset, exec_instr{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}
	cp_cfg_A_na4_r : cross legal_RWX_L_NA4, addr_offset, read_instr_lw{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}
	cp_cfg_A_na4_w : cross legal_RWX_L_NA4, addr_offset, write_instr_sw{
		ignore_bins ig1  = binsof(addr_offset.below_base);
		ignore_bins ig2  = binsof(addr_offset.highest_word);
	}

	cp_cfg_A_NA4_all: cross pmpcfgA_NA4, RWXL001, read_instr_lw, addr_offset{
		ignore_bins ig5  = binsof(addr_offset.just_beyond);
		ignore_bins ig6  = binsof(addr_offset.highest_word);
	}

	cp_pmpaddr_walk: cross priv_mode_m, cp_walk_rs1_pmpaddr, csrrw, legal_pmpaddr_entries ;
	cp_pmpcfg_walk: cross priv_mode_m, cp_walk_rs1_pmpcfg, csrrw, legal_pmpcfg_entries_even ;
	cp_pmpcfg_zero: cross priv_mode_m, cp_zero_rs1, csrrw, legal_pmpcfg_entries_odd ;

	cp_pmp64_write: cross priv_mode_m, write_instr_sw, pmp64;
	cp_pmp64_read: cross priv_mode_m, read_instr_lw, pmp64;

endgroup

function void pmp_sample(int hart, int issue, ins_t ins);

	logic [XLEN-1:0] pmpcfg [15:0];
	logic [XLEN-1:0] pmpaddr [62:0];
	logic [29:0] pmpcfg_rw, pmpcfg_a;			// for first 15 Regions
	logic [95:0] pmpcfg_RW, pmpcfg_A;			// for next 48 Regions
	logic [14:0] pmpcfg_x, pmpcfg_l, pmp_hit;   // for first 15 Regions
	logic [47:0] pmpcfg_X, pmpcfg_L, pmp_HIT;   // for next 48 Regions

	for (int i = 0; i < 16; i++) begin
		pmpcfg[i] = ins.current.csr[12'h3A0 + i];
	end

	for (int j = 0; j < 63; j++) begin
		pmpaddr[j] = ins.current.csr[12'h3B0 + j];
	end

	for (int k = 0; k < 15; k++) begin				// for first 15 regions
		pmp_hit[k] = (pmpaddr[k] == `REGIONSTART);
	end

	for (int k = 15; k < 64; k++) begin				// for next 48 regions
		pmp_HIT[k] = (pmpaddr[k] == `REGIONSTART);
	end

	`ifdef XLEN32
		pmpcfg_rw = {
					ins.current.csr[12'h3A3][17:16],
					ins.current.csr[12'h3A3][9:8],
					ins.current.csr[12'h3A3][1:0],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A1][25:24],
					ins.current.csr[12'h3A1][17:16],
					ins.current.csr[12'h3A1][9:8],
					ins.current.csr[12'h3A1][1:0],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_rw = {
					ins.current.csr[12'h3A2][49:48],
					ins.current.csr[12'h3A2][41:40],
					ins.current.csr[12'h3A2][33:32],
					ins.current.csr[12'h3A2][25:24],
					ins.current.csr[12'h3A2][17:16],
					ins.current.csr[12'h3A2][9:8],
					ins.current.csr[12'h3A2][1:0],
					ins.current.csr[12'h3A0][57:56],
					ins.current.csr[12'h3A0][49:48],
					ins.current.csr[12'h3A0][41:40],
					ins.current.csr[12'h3A0][33:32],
					ins.current.csr[12'h3A0][25:24],
					ins.current.csr[12'h3A0][17:16],
					ins.current.csr[12'h3A0][9:8],
					ins.current.csr[12'h3A0][1:0]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_RW = {
					ins.current.csr[12'h3AF][17:16],
					ins.current.csr[12'h3AF][9:8],
					ins.current.csr[12'h3AF][1:0],
					ins.current.csr[12'h3AE][25:24],
					ins.current.csr[12'h3AE][17:16],
					ins.current.csr[12'h3AE][9:8],
					ins.current.csr[12'h3AE][1:0],
					ins.current.csr[12'h3AD][25:24],
					ins.current.csr[12'h3AD][17:16],
					ins.current.csr[12'h3AD][9:8],
					ins.current.csr[12'h3AD][1:0],
					ins.current.csr[12'h3AC][25:24],
					ins.current.csr[12'h3AC][17:16],
					ins.current.csr[12'h3AC][9:8],
					ins.current.csr[12'h3AC][1:0],
					ins.current.csr[12'h3AB][25:24],
					ins.current.csr[12'h3AB][17:16],
					ins.current.csr[12'h3AB][9:8],
					ins.current.csr[12'h3AB][1:0],
					ins.current.csr[12'h3AA][25:24],
					ins.current.csr[12'h3AA][17:16],
					ins.current.csr[12'h3AA][9:8],
					ins.current.csr[12'h3AA][1:0],
					ins.current.csr[12'h3A9][25:24],
					ins.current.csr[12'h3A9][17:16],
					ins.current.csr[12'h3A9][9:8],
					ins.current.csr[12'h3A9][1:0],
					ins.current.csr[12'h3A8][25:24],
					ins.current.csr[12'h3A8][17:16],
					ins.current.csr[12'h3A8][9:8],
					ins.current.csr[12'h3A8][1:0],
					ins.current.csr[12'h3A7][25:24],
					ins.current.csr[12'h3A7][17:16],
					ins.current.csr[12'h3A7][9:8],
					ins.current.csr[12'h3A7][1:0],
					ins.current.csr[12'h3A6][25:24],
					ins.current.csr[12'h3A6][17:16],
					ins.current.csr[12'h3A6][9:8],
					ins.current.csr[12'h3A6][1:0],
					ins.current.csr[12'h3A5][25:24],
					ins.current.csr[12'h3A5][17:16],
					ins.current.csr[12'h3A5][9:8],
					ins.current.csr[12'h3A5][1:0],
					ins.current.csr[12'h3A4][25:24],
					ins.current.csr[12'h3A4][17:16],
					ins.current.csr[12'h3A4][9:8],
					ins.current.csr[12'h3A4][1:0],
					ins.current.csr[12'h3A3][25:24]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_RW = {
					ins.current.csr[12'h3AE][49:48],
					ins.current.csr[12'h3AE][41:40],
					ins.current.csr[12'h3AE][33:32],
					ins.current.csr[12'h3AE][25:24],
					ins.current.csr[12'h3AE][17:16],
					ins.current.csr[12'h3AE][9:8],
					ins.current.csr[12'h3AE][1:0],
					ins.current.csr[12'h3AC][57:56],
					ins.current.csr[12'h3AC][49:48],
					ins.current.csr[12'h3AC][41:40],
					ins.current.csr[12'h3AC][33:32],
					ins.current.csr[12'h3AC][25:24],
					ins.current.csr[12'h3AC][17:16],
					ins.current.csr[12'h3AC][9:8],
					ins.current.csr[12'h3AC][1:0],
					ins.current.csr[12'h3AA][57:56],
					ins.current.csr[12'h3AA][49:48],
					ins.current.csr[12'h3AA][41:40],
					ins.current.csr[12'h3AA][33:32],
					ins.current.csr[12'h3AA][25:24],
					ins.current.csr[12'h3AA][17:16],
					ins.current.csr[12'h3AA][9:8],
					ins.current.csr[12'h3AA][1:0],
					ins.current.csr[12'h3A8][57:56],
					ins.current.csr[12'h3A8][49:48],
					ins.current.csr[12'h3A8][41:40],
					ins.current.csr[12'h3A8][33:32],
					ins.current.csr[12'h3A8][25:24],
					ins.current.csr[12'h3A8][17:16],
					ins.current.csr[12'h3A8][9:8],
					ins.current.csr[12'h3A8][1:0],
					ins.current.csr[12'h3A6][57:56],
					ins.current.csr[12'h3A6][49:48],
					ins.current.csr[12'h3A6][41:40],
					ins.current.csr[12'h3A6][33:32],
					ins.current.csr[12'h3A6][25:24],
					ins.current.csr[12'h3A6][17:16],
					ins.current.csr[12'h3A6][9:8],
					ins.current.csr[12'h3A6][1:0],
					ins.current.csr[12'h3A4][57:56],
					ins.current.csr[12'h3A4][49:48],
					ins.current.csr[12'h3A4][41:40],
					ins.current.csr[12'h3A4][33:32],
					ins.current.csr[12'h3A4][25:24],
					ins.current.csr[12'h3A4][17:16],
					ins.current.csr[12'h3A4][9:8],
					ins.current.csr[12'h3A4][1:0],
					ins.current.csr[12'h3A2][57:56]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_X =  {
					ins.current.csr[12'h3AF][18],
					ins.current.csr[12'h3AF][10],
					ins.current.csr[12'h3AF][2],
					ins.current.csr[12'h3AE][26],
					ins.current.csr[12'h3AE][18],
					ins.current.csr[12'h3AE][10],
					ins.current.csr[12'h3AE][2],
					ins.current.csr[12'h3AD][26],
					ins.current.csr[12'h3AD][18],
					ins.current.csr[12'h3AD][10],
					ins.current.csr[12'h3AD][2],
					ins.current.csr[12'h3AC][26],
					ins.current.csr[12'h3AC][18],
					ins.current.csr[12'h3AC][10],
					ins.current.csr[12'h3AC][2],
					ins.current.csr[12'h3AB][26],
					ins.current.csr[12'h3AB][18],
					ins.current.csr[12'h3AB][10],
					ins.current.csr[12'h3AB][2],
					ins.current.csr[12'h3AA][26],
					ins.current.csr[12'h3AA][18],
					ins.current.csr[12'h3AA][10],
					ins.current.csr[12'h3AA][2],
					ins.current.csr[12'h3A9][26],
					ins.current.csr[12'h3A9][18],
					ins.current.csr[12'h3A9][10],
					ins.current.csr[12'h3A9][2],
					ins.current.csr[12'h3A8][26],
					ins.current.csr[12'h3A8][18],
					ins.current.csr[12'h3A8][10],
					ins.current.csr[12'h3A8][2],
					ins.current.csr[12'h3A7][26],
					ins.current.csr[12'h3A7][18],
					ins.current.csr[12'h3A7][10],
					ins.current.csr[12'h3A7][2],
					ins.current.csr[12'h3A6][26],
					ins.current.csr[12'h3A6][18],
					ins.current.csr[12'h3A6][10],
					ins.current.csr[12'h3A6][2],
					ins.current.csr[12'h3A5][26],
					ins.current.csr[12'h3A5][18],
					ins.current.csr[12'h3A5][10],
					ins.current.csr[12'h3A5][2],
					ins.current.csr[12'h3A4][26],
					ins.current.csr[12'h3A4][18],
					ins.current.csr[12'h3A4][10],
					ins.current.csr[12'h3A4][2],
					ins.current.csr[12'h3A3][18]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_X =  {
					ins.current.csr[12'h3AE][50],
					ins.current.csr[12'h3AE][42],
					ins.current.csr[12'h3AE][34],
					ins.current.csr[12'h3AE][26],
					ins.current.csr[12'h3AE][18],
					ins.current.csr[12'h3AE][10],
					ins.current.csr[12'h3AE][2],
					ins.current.csr[12'h3AC][58],
					ins.current.csr[12'h3AC][50],
					ins.current.csr[12'h3AC][42],
					ins.current.csr[12'h3AC][34],
					ins.current.csr[12'h3AC][26],
					ins.current.csr[12'h3AC][18],
					ins.current.csr[12'h3AC][10],
					ins.current.csr[12'h3AC][2],
					ins.current.csr[12'h3AA][58],
					ins.current.csr[12'h3AA][50],
					ins.current.csr[12'h3AA][42],
					ins.current.csr[12'h3AA][34],
					ins.current.csr[12'h3AA][26],
					ins.current.csr[12'h3AA][18],
					ins.current.csr[12'h3AA][10],
					ins.current.csr[12'h3AA][2],
					ins.current.csr[12'h3A8][58],
					ins.current.csr[12'h3A8][50],
					ins.current.csr[12'h3A8][42],
					ins.current.csr[12'h3A8][34],
					ins.current.csr[12'h3A8][26],
					ins.current.csr[12'h3A8][18],
					ins.current.csr[12'h3A8][10],
					ins.current.csr[12'h3A8][2],
					ins.current.csr[12'h3A6][58],
					ins.current.csr[12'h3A6][50],
					ins.current.csr[12'h3A6][42],
					ins.current.csr[12'h3A6][34],
					ins.current.csr[12'h3A6][26],
					ins.current.csr[12'h3A6][18],
					ins.current.csr[12'h3A6][10],
					ins.current.csr[12'h3A6][2],
					ins.current.csr[12'h3A4][58],
					ins.current.csr[12'h3A4][50],
					ins.current.csr[12'h3A4][42],
					ins.current.csr[12'h3A4][34],
					ins.current.csr[12'h3A4][26],
					ins.current.csr[12'h3A4][18],
					ins.current.csr[12'h3A4][10],
					ins.current.csr[12'h3A4][2],
					ins.current.csr[12'h3A2][58]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_x =  {
					ins.current.csr[12'h3A3][18],
					ins.current.csr[12'h3A3][10],
					ins.current.csr[12'h3A3][2],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A1][26],
					ins.current.csr[12'h3A1][18],
					ins.current.csr[12'h3A1][10],
					ins.current.csr[12'h3A1][2],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_x =  {
					ins.current.csr[12'h3A2][50],
					ins.current.csr[12'h3A2][42],
					ins.current.csr[12'h3A2][34],
					ins.current.csr[12'h3A2][26],
					ins.current.csr[12'h3A2][18],
					ins.current.csr[12'h3A2][10],
					ins.current.csr[12'h3A2][2],
					ins.current.csr[12'h3A0][58],
					ins.current.csr[12'h3A0][50],
					ins.current.csr[12'h3A0][42],
					ins.current.csr[12'h3A0][34],
					ins.current.csr[12'h3A0][26],
					ins.current.csr[12'h3A0][18],
					ins.current.csr[12'h3A0][10],
					ins.current.csr[12'h3A0][2]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_a =  {
					ins.current.csr[12'h3A3][20:19],
					ins.current.csr[12'h3A3][12:11],
					ins.current.csr[12'h3A3][4:3],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A1][28:27],
					ins.current.csr[12'h3A1][20:19],
					ins.current.csr[12'h3A1][12:11],
					ins.current.csr[12'h3A1][4:3],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_a =  {
					ins.current.csr[12'h3A2][52:51],
					ins.current.csr[12'h3A2][44:43],
					ins.current.csr[12'h3A2][36:35],
					ins.current.csr[12'h3A2][28:27],
					ins.current.csr[12'h3A2][20:19],
					ins.current.csr[12'h3A2][12:11],
					ins.current.csr[12'h3A2][4:3],
					ins.current.csr[12'h3A0][60:59],
					ins.current.csr[12'h3A0][52:51],
					ins.current.csr[12'h3A0][44:43],
					ins.current.csr[12'h3A0][36:35],
					ins.current.csr[12'h3A0][28:27],
					ins.current.csr[12'h3A0][20:19],
					ins.current.csr[12'h3A0][12:11],
					ins.current.csr[12'h3A0][4:3]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_A =  {
					ins.current.csr[12'h3AF][20:19],
					ins.current.csr[12'h3AF][12:11],
					ins.current.csr[12'h3AF][4:3],
					ins.current.csr[12'h3AE][28:27],
					ins.current.csr[12'h3AE][20:19],
					ins.current.csr[12'h3AE][12:11],
					ins.current.csr[12'h3AE][4:3],
					ins.current.csr[12'h3AD][28:27],
					ins.current.csr[12'h3AD][20:19],
					ins.current.csr[12'h3AD][12:11],
					ins.current.csr[12'h3AD][4:3],
					ins.current.csr[12'h3AC][28:27],
					ins.current.csr[12'h3AC][20:19],
					ins.current.csr[12'h3AC][12:11],
					ins.current.csr[12'h3AC][4:3],
					ins.current.csr[12'h3AB][28:27],
					ins.current.csr[12'h3AB][20:19],
					ins.current.csr[12'h3AB][12:11],
					ins.current.csr[12'h3AB][4:3],
					ins.current.csr[12'h3AA][28:27],
					ins.current.csr[12'h3AA][20:19],
					ins.current.csr[12'h3AA][12:11],
					ins.current.csr[12'h3AA][4:3],
					ins.current.csr[12'h3A9][28:27],
					ins.current.csr[12'h3A9][20:19],
					ins.current.csr[12'h3A9][12:11],
					ins.current.csr[12'h3A9][4:3],
					ins.current.csr[12'h3A8][28:27],
					ins.current.csr[12'h3A8][20:19],
					ins.current.csr[12'h3A8][12:11],
					ins.current.csr[12'h3A8][4:3],
					ins.current.csr[12'h3A7][28:27],
					ins.current.csr[12'h3A7][20:19],
					ins.current.csr[12'h3A7][12:11],
					ins.current.csr[12'h3A7][4:3],
					ins.current.csr[12'h3A6][28:27],
					ins.current.csr[12'h3A6][20:19],
					ins.current.csr[12'h3A6][12:11],
					ins.current.csr[12'h3A6][4:3],
					ins.current.csr[12'h3A5][28:27],
					ins.current.csr[12'h3A5][20:19],
					ins.current.csr[12'h3A5][12:11],
					ins.current.csr[12'h3A5][4:3],
					ins.current.csr[12'h3A4][28:27],
					ins.current.csr[12'h3A4][20:19],
					ins.current.csr[12'h3A4][12:11],
					ins.current.csr[12'h3A4][4:3],
					ins.current.csr[12'h3A3][28:27]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_A =  {
					ins.current.csr[12'h3AE][52:51],
					ins.current.csr[12'h3AE][44:43],
					ins.current.csr[12'h3AE][36:35],
					ins.current.csr[12'h3AE][28:27],
					ins.current.csr[12'h3AE][20:19],
					ins.current.csr[12'h3AE][12:11],
					ins.current.csr[12'h3AE][4:3],
					ins.current.csr[12'h3AC][60:59],
					ins.current.csr[12'h3AC][52:51],
					ins.current.csr[12'h3AC][44:43],
					ins.current.csr[12'h3AC][36:35],
					ins.current.csr[12'h3AC][28:27],
					ins.current.csr[12'h3AC][20:19],
					ins.current.csr[12'h3AC][12:11],
					ins.current.csr[12'h3AC][4:3],
					ins.current.csr[12'h3AA][60:59],
					ins.current.csr[12'h3AA][52:51],
					ins.current.csr[12'h3AA][44:43],
					ins.current.csr[12'h3AA][36:35],
					ins.current.csr[12'h3AA][28:27],
					ins.current.csr[12'h3AA][20:19],
					ins.current.csr[12'h3AA][12:11],
					ins.current.csr[12'h3AA][4:3],
					ins.current.csr[12'h3A8][60:59],
					ins.current.csr[12'h3A8][52:51],
					ins.current.csr[12'h3A8][44:43],
					ins.current.csr[12'h3A8][36:35],
					ins.current.csr[12'h3A8][28:27],
					ins.current.csr[12'h3A8][20:19],
					ins.current.csr[12'h3A8][12:11],
					ins.current.csr[12'h3A8][4:3],
					ins.current.csr[12'h3A6][60:59],
					ins.current.csr[12'h3A6][52:51],
					ins.current.csr[12'h3A6][44:43],
					ins.current.csr[12'h3A6][36:35],
					ins.current.csr[12'h3A6][28:27],
					ins.current.csr[12'h3A6][20:19],
					ins.current.csr[12'h3A6][12:11],
					ins.current.csr[12'h3A6][4:3],
					ins.current.csr[12'h3A4][60:59],
					ins.current.csr[12'h3A4][52:51],
					ins.current.csr[12'h3A4][44:43],
					ins.current.csr[12'h3A4][36:35],
					ins.current.csr[12'h3A4][28:27],
					ins.current.csr[12'h3A4][20:19],
					ins.current.csr[12'h3A4][12:11],
					ins.current.csr[12'h3A4][4:3],
					ins.current.csr[12'h3A2][60:59]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_L =  {
					ins.current.csr[12'h3AF][23],
					ins.current.csr[12'h3AF][15],
					ins.current.csr[12'h3AF][7],
					ins.current.csr[12'h3AD][31],
					ins.current.csr[12'h3AD][23],
					ins.current.csr[12'h3AD][15],
					ins.current.csr[12'h3AD][7],
					ins.current.csr[12'h3AD][31],
					ins.current.csr[12'h3AD][23],
					ins.current.csr[12'h3AD][15],
					ins.current.csr[12'h3AD][7],
					ins.current.csr[12'h3AC][31],
					ins.current.csr[12'h3AC][23],
					ins.current.csr[12'h3AC][15],
					ins.current.csr[12'h3AC][7],
					ins.current.csr[12'h3AB][31],
					ins.current.csr[12'h3AB][23],
					ins.current.csr[12'h3AB][15],
					ins.current.csr[12'h3AB][7],
					ins.current.csr[12'h3AA][31],
					ins.current.csr[12'h3AA][23],
					ins.current.csr[12'h3AA][15],
					ins.current.csr[12'h3AA][7],
					ins.current.csr[12'h3A9][31],
					ins.current.csr[12'h3A9][23],
					ins.current.csr[12'h3A9][15],
					ins.current.csr[12'h3A9][7],
					ins.current.csr[12'h3A8][31],
					ins.current.csr[12'h3A8][23],
					ins.current.csr[12'h3A8][15],
					ins.current.csr[12'h3A8][7],
					ins.current.csr[12'h3A7][31],
					ins.current.csr[12'h3A7][23],
					ins.current.csr[12'h3A7][15],
					ins.current.csr[12'h3A7][7],
					ins.current.csr[12'h3A6][31],
					ins.current.csr[12'h3A6][23],
					ins.current.csr[12'h3A6][15],
					ins.current.csr[12'h3A6][7],
					ins.current.csr[12'h3A5][31],
					ins.current.csr[12'h3A5][23],
					ins.current.csr[12'h3A5][15],
					ins.current.csr[12'h3A5][7],
					ins.current.csr[12'h3A4][31],
					ins.current.csr[12'h3A4][23],
					ins.current.csr[12'h3A4][15],
					ins.current.csr[12'h3A4][7],
					ins.current.csr[12'h3A3][31]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_L =  {
					ins.current.csr[12'h3AE][55],
					ins.current.csr[12'h3AE][47],
					ins.current.csr[12'h3AE][39],
					ins.current.csr[12'h3AE][31],
					ins.current.csr[12'h3AE][23],
					ins.current.csr[12'h3AE][15],
					ins.current.csr[12'h3AE][7],
					ins.current.csr[12'h3AC][63],
					ins.current.csr[12'h3AC][55],
					ins.current.csr[12'h3AC][47],
					ins.current.csr[12'h3AC][39],
					ins.current.csr[12'h3AC][31],
					ins.current.csr[12'h3AC][23],
					ins.current.csr[12'h3AC][15],
					ins.current.csr[12'h3AC][7],
					ins.current.csr[12'h3AA][63]
					ins.current.csr[12'h3AA][55],
					ins.current.csr[12'h3AA][47],
					ins.current.csr[12'h3AA][39],
					ins.current.csr[12'h3AA][31],
					ins.current.csr[12'h3AA][23],
					ins.current.csr[12'h3AA][15],
					ins.current.csr[12'h3AA][7],
					ins.current.csr[12'h3A8][63],
					ins.current.csr[12'h3A8][55],
					ins.current.csr[12'h3A8][47],
					ins.current.csr[12'h3A8][39],
					ins.current.csr[12'h3A8][31],
					ins.current.csr[12'h3A8][23],
					ins.current.csr[12'h3A8][15],
					ins.current.csr[12'h3A8][7],
					ins.current.csr[12'h3A6][63]
					ins.current.csr[12'h3A6][55],
					ins.current.csr[12'h3A6][47],
					ins.current.csr[12'h3A6][39],
					ins.current.csr[12'h3A6][31],
					ins.current.csr[12'h3A6][23],
					ins.current.csr[12'h3A6][15],
					ins.current.csr[12'h3A6][7],
					ins.current.csr[12'h3A4][63],
					ins.current.csr[12'h3A4][55],
					ins.current.csr[12'h3A4][47],
					ins.current.csr[12'h3A4][39],
					ins.current.csr[12'h3A4][31],
					ins.current.csr[12'h3A4][23],
					ins.current.csr[12'h3A4][15],
					ins.current.csr[12'h3A4][7],
					ins.current.csr[12'h3A2][63]
					};
	`endif

	`ifdef XLEN32
		pmpcfg_l =  {
					ins.current.csr[12'h3A3][23],
					ins.current.csr[12'h3A3][15],
					ins.current.csr[12'h3A3][7],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A1][31],
					ins.current.csr[12'h3A1][23],
					ins.current.csr[12'h3A1][15],
					ins.current.csr[12'h3A1][7],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif
	`ifdef XLEN64
		pmpcfg_l =  {
					ins.current.csr[12'h3A2][55],
					ins.current.csr[12'h3A2][47],
					ins.current.csr[12'h3A2][39],
					ins.current.csr[12'h3A2][31],
					ins.current.csr[12'h3A2][23],
					ins.current.csr[12'h3A2][15],
					ins.current.csr[12'h3A2][7],
					ins.current.csr[12'h3A0][63],
					ins.current.csr[12'h3A0][55],
					ins.current.csr[12'h3A0][47],
					ins.current.csr[12'h3A0][39],
					ins.current.csr[12'h3A0][31],
					ins.current.csr[12'h3A0][23],
					ins.current.csr[12'h3A0][15],
					ins.current.csr[12'h3A0][7]
					};
	`endif

	PMPM_cg.sample(ins, pmpcfg, pmpaddr, pmpcfg_rw, pmpcfg_RW, pmpcfg_a, pmpcfg_A, pmpcfg_x, pmpcfg_X, pmpcfg_l, pmpcfg_L, pmp_hit, pmp_HIT);
endfunction
