///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    csrrc_cg = new(); csrrc_cg.set_inst_name("obj_csrrc");
    csrrci_cg = new(); csrrci_cg.set_inst_name("obj_csrrci");
    csrrs_cg = new(); csrrs_cg.set_inst_name("obj_csrrs");
    csrrsi_cg = new(); csrrsi_cg.set_inst_name("obj_csrrsi");
    csrrw_cg = new(); csrrw_cg.set_inst_name("obj_csrrw");
    csrrwi_cg = new(); csrrwi_cg.set_inst_name("obj_csrrwi");
