///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    andn_cg = new(); andn_cg.set_inst_name("obj_andn");
    clz_cg = new(); clz_cg.set_inst_name("obj_clz");
    clzw_cg = new(); clzw_cg.set_inst_name("obj_clzw");
    cpop_cg = new(); cpop_cg.set_inst_name("obj_cpop");
    cpopw_cg = new(); cpopw_cg.set_inst_name("obj_cpopw");
    ctz_cg = new(); ctz_cg.set_inst_name("obj_ctz");
    ctzw_cg = new(); ctzw_cg.set_inst_name("obj_ctzw");
    max_cg = new(); max_cg.set_inst_name("obj_max");
    maxu_cg = new(); maxu_cg.set_inst_name("obj_maxu");
    min_cg = new(); min_cg.set_inst_name("obj_min");
    minu_cg = new(); minu_cg.set_inst_name("obj_minu");
    orc_b_cg = new(); orc_b_cg.set_inst_name("obj_orc_b");
    orn_cg = new(); orn_cg.set_inst_name("obj_orn");
    rev8_cg = new(); rev8_cg.set_inst_name("obj_rev8");
    rol_cg = new(); rol_cg.set_inst_name("obj_rol");
    rolw_cg = new(); rolw_cg.set_inst_name("obj_rolw");
    ror_cg = new(); ror_cg.set_inst_name("obj_ror");
    rori_cg = new(); rori_cg.set_inst_name("obj_rori");
    roriw_cg = new(); roriw_cg.set_inst_name("obj_roriw");
    rorw_cg = new(); rorw_cg.set_inst_name("obj_rorw");
    sext_b_cg = new(); sext_b_cg.set_inst_name("obj_sext_b");
    sext_h_cg = new(); sext_h_cg.set_inst_name("obj_sext_h");
    xnor_cg = new(); xnor_cg.set_inst_name("obj_xnor");
    zext_h_cg = new(); zext_h_cg.set_inst_name("obj_zext_h");
