///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    fadd_h_cg = new(); fadd_h_cg.set_inst_name("obj_fadd_h");
    fclass_h_cg = new(); fclass_h_cg.set_inst_name("obj_fclass_h");
    fcvt_h_s_cg = new(); fcvt_h_s_cg.set_inst_name("obj_fcvt_h_s");
    fcvt_h_w_cg = new(); fcvt_h_w_cg.set_inst_name("obj_fcvt_h_w");
    fcvt_h_wu_cg = new(); fcvt_h_wu_cg.set_inst_name("obj_fcvt_h_wu");
    fcvt_s_h_cg = new(); fcvt_s_h_cg.set_inst_name("obj_fcvt_s_h");
    fcvt_w_h_cg = new(); fcvt_w_h_cg.set_inst_name("obj_fcvt_w_h");
    fcvt_wu_h_cg = new(); fcvt_wu_h_cg.set_inst_name("obj_fcvt_wu_h");
    fdiv_h_cg = new(); fdiv_h_cg.set_inst_name("obj_fdiv_h");
    feq_h_cg = new(); feq_h_cg.set_inst_name("obj_feq_h");
    fle_h_cg = new(); fle_h_cg.set_inst_name("obj_fle_h");
    flh_cg = new(); flh_cg.set_inst_name("obj_flh");
    flt_h_cg = new(); flt_h_cg.set_inst_name("obj_flt_h");
    fmadd_h_cg = new(); fmadd_h_cg.set_inst_name("obj_fmadd_h");
    fmax_h_cg = new(); fmax_h_cg.set_inst_name("obj_fmax_h");
    fmin_h_cg = new(); fmin_h_cg.set_inst_name("obj_fmin_h");
    fmsub_h_cg = new(); fmsub_h_cg.set_inst_name("obj_fmsub_h");
    fmul_h_cg = new(); fmul_h_cg.set_inst_name("obj_fmul_h");
    fmv_h_x_cg = new(); fmv_h_x_cg.set_inst_name("obj_fmv_h_x");
    fmv_x_h_cg = new(); fmv_x_h_cg.set_inst_name("obj_fmv_x_h");
    fnmadd_h_cg = new(); fnmadd_h_cg.set_inst_name("obj_fnmadd_h");
    fnmsub_h_cg = new(); fnmsub_h_cg.set_inst_name("obj_fnmsub_h");
    fsgnj_h_cg = new(); fsgnj_h_cg.set_inst_name("obj_fsgnj_h");
    fsgnjn_h_cg = new(); fsgnjn_h_cg.set_inst_name("obj_fsgnjn_h");
    fsgnjx_h_cg = new(); fsgnjx_h_cg.set_inst_name("obj_fsgnjx_h");
    fsh_cg = new(); fsh_cg.set_inst_name("obj_fsh");
    fsqrt_h_cg = new(); fsqrt_h_cg.set_inst_name("obj_fsqrt_h");
    fsub_h_cg = new(); fsub_h_cg.set_inst_name("obj_fsub_h");
