///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ExceptionsV_edgecases_cg = new();           ExceptionsV_edgecases_cg.set_inst_name("obj_ExceptionsV_edgecases");
    ExceptionsV_reserved_cg = new();            ExceptionsV_reserved_cg.set_inst_name("obj_ExceptionsV_reserved");
    ExceptionsV_illegal_cg = new();             ExceptionsV_illegal_cg.set_inst_name("obj_ExceptionsV_illegal");
