///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    aes32esi_cg = new(); aes32esi_cg.set_inst_name("obj_aes32esi");
    aes32esmi_cg = new(); aes32esmi_cg.set_inst_name("obj_aes32esmi");
