///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    scsr_cg = new();        scsr_cg.set_inst_name("obj_scsr");
    scause_cg = new();      scause_cg.set_inst_name("obj_scause");
    sstatus_cg = new();     sstatus_cg.set_inst_name("obj_sstatus");
    sprivinst_cg = new();   sprivinst_cg.set_inst_name("obj_sprivinst");

 
