///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    andn_cg = new(); andn_cg.set_inst_name("obj_andn");
    brev8_cg = new(); brev8_cg.set_inst_name("obj_brev8");
    orn_cg = new(); orn_cg.set_inst_name("obj_orn");
    pack_cg = new(); pack_cg.set_inst_name("obj_pack");
    packh_cg = new(); packh_cg.set_inst_name("obj_packh");
    rev8_cg = new(); rev8_cg.set_inst_name("obj_rev8");
    rol_cg = new(); rol_cg.set_inst_name("obj_rol");
    ror_cg = new(); ror_cg.set_inst_name("obj_ror");
    rori_cg = new(); rori_cg.set_inst_name("obj_rori");
    xor_cg = new(); xor_cg.set_inst_name("obj_xor");
