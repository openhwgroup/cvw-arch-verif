///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Written: Corey Hickson chickson@hmc.edu, Jordan Carlin jcarlin@hmc.edu 08 Feb 2025
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_INTERRUPTSM
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_interruptsm_t;

covergroup InterruptsM_cg with function sample(ins_interruptsm_t ins);
    option.per_instance = 0; 

    // building blocks for the main coverpoints
    
    mstatus_mie_one: coverpoint ins.current.csr[12'h300][3] {
        bins zero = {1};
    }
    mstatus_mie: coverpoint ins.current.csr[12'h300][3]  {
        // autofill 0/1
    }
    mstatus_tw:  coverpoint ins.current.csr[12'h300][21] {
        // autofill 0/1
    }

    mie_mtie_one: coverpoint ins.current.csr[12'h304][7] {
        bins one = {1};
    }
    mie_ones: coverpoint ins.current.csr[12'h304][15:0] {
        wildcard bins ones = {16'b????1???1???1???}; // ones in every field that is not tied to zero
    }
    mip_msip_one: coverpoint ins.current.csr[12'h344][3] {
        bins one = {1};
    }
    mip_mtip: coverpoint ins.current.csr[12'h344][7] {
        // autofill 0/1
    }
    mip_mtip_one: coverpoint ins.current.csr[12'h344][7] {
        bins one = {1};
    }
    mip_meip_one: coverpoint ins.current.csr[12'h344][11] {
        bins one = {1};
    }
    mie_walking: coverpoint {ins.current.csr[12'h304][11],
                             ins.current.csr[12'h304][7], 
                             ins.current.csr[12'h304][3] } {
        bins meie = {3'b001};
        bins mtie = {3'b010};
        bins msie = {3'b100};
    }
    mip_walking: coverpoint {ins.current.csr[12'h344][11],
                             ins.current.csr[12'h344][7], 
                             ins.current.csr[12'h344][3] } {
        bins meip = {3'b001};
        bins mtip = {3'b010};
        bins msip = {3'b100};
    }
    mie_meie_mtie_msie: coverpoint {ins.current.csr[12'h304][11],
                                    ins.current.csr[12'h304][7], 
                                    ins.current.csr[12'h304][3] } {
        // auto fills all 8 combinations
    }
    mip_meip_mtip_msip: coverpoint {ins.current.csr[12'h344][11],
                                    ins.current.csr[12'h344][7], 
                                    ins.current.csr[12'h344][3] } {
        // auto fills all 8 combinations
    }
    mtvec_direct: coverpoint ins.current.csr[12'h305][1:0] {
        bins direct   = {2'b00};
    }
    mtvec_vectored: coverpoint ins.current.csr[12'h305][1:0] {
        bins vector   = {2'b01};
    }
    wfi: coverpoint ins.current.insn {
        bins wfi = {32'b0001000_00101_00000_000_00000_1110011};
    }
    priv_mode_m: coverpoint ins.current.mode {
        bins M_mode = {2'b11};
    }
    m_ext_intr: coverpoint ins.current.m_ext_intr {
        bins mei = {1};
    }
    m_timer_intr: coverpoint ins.current.m_timer_intr {
        bins mti = {1};
    }
    m_soft_intr: coverpoint ins.current.m_soft_intr {
        bins msi = {1};
    }

    // main coverpoints

    cp_trigger_mti:      cross priv_mode_m, mstatus_mie, mie_ones, m_timer_intr, mip_mtip_one; // redundant to check both?
    cp_trigger_msi:      cross priv_mode_m, mstatus_mie, mie_ones, m_soft_intr,  mip_msip_one; // if not, should we check rising
    cp_trigger_mei:      cross priv_mode_m, mstatus_mie, mie_ones, m_ext_intr,   mip_meip_one; // edge transitions for m*ip?
    cp_global_ie:        cross priv_mode_m, mstatus_mie, mip_walking, mie_walking;
    cp_interrupts:       cross priv_mode_m, mstatus_mie, mtvec_direct, mip_walking, mie_walking;
    cp_vectored:         cross priv_mode_m, mstatus_mie_one, mtvec_vectored, mip_walking, mie_walking;
    cp_priority:         cross priv_mode_m, mstatus_mie_one, mie_meie_mtie_msie, mip_meip_mtip_msip;
    cp_wfi:              cross priv_mode_m, wfi, mstatus_mie, mstatus_tw, mie_mtie_one, m_timer_intr;
endgroup

function void interruptsm_sample(int hart, int issue);
    ins_interruptsm_t ins;

    ins = new(hart, issue, traceDataQ); 
    ins.add_rd(0);
    ins.add_rs1(2);
    ins.add_csr(1);
    
    InterruptsM_cg.sample(ins);
    
endfunction
