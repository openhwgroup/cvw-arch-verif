///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    SsstrictS_instr_cg = new();        SsstrictS_instr_cg.set_inst_name("obj_SsstrictS_instr");
    SsstrictS_comp_instr_cg = new();   SsstrictS_comp_instr_cg.set_inst_name("obj_SsstrictS_comp_instr");
    SsstrictS_scsr_cg = new();         SsstrictS_scsr_cg.set_inst_name("obj_SsstrictS_scsr");
     
