///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    xperm4_cg = new(); xperm4_cg.set_inst_name("obj_xperm4");
    xperm8_cg = new(); xperm8_cg.set_inst_name("obj_xperm8");
