///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_RV64I
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_rv64i_t;


covergroup add_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "add";
    cp_asm_count : coverpoint ins.ins_str == "add"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup addi_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "addi";
    cp_asm_count : coverpoint ins.ins_str == "addi"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup addiw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "addiw";
    cp_asm_count : coverpoint ins.ins_str == "addiw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup addw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "addw";
    cp_asm_count : coverpoint ins.ins_str == "addw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup and_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "and";
    cp_asm_count : coverpoint ins.ins_str == "and"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup andi_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "andi";
    cp_asm_count : coverpoint ins.ins_str == "andi"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup auipc_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "auipc";
    cp_asm_count : coverpoint ins.ins_str == "auipc"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle_auipc : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners for auipc";
        wildcard bins bit_12_0 = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0 = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0 = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0 = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0 = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0 = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0 = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0 = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0 = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0 = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0 = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0 = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0 = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0 = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0 = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0 = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0 = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0 = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0 = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0 = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0 = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0 = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0 = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0 = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0 = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0 = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0 = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0 = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0 = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0 = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0 = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0 = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0 = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0 = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0 = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0 = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0 = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0 = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0 = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0 = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0 = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0 = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0 = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0 = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0 = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0 = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0 = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0 = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0 = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0 = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0 = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0 = {64'b0???????????????????????????????????????????????????????????????};

        wildcard bins bit_12_1 = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1 = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1 = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1 = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1 = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1 = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1 = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1 = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1 = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1 = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1 = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1 = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1 = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1 = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1 = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1 = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1 = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1 = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1 = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1 = {64'b????????????????????????????????1???????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm_zero : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        bins zero  = {0};
        bins nonzero  = default;
    }
endgroup

covergroup beq_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "beq";
    cp_asm_count : coverpoint ins.ins_str == "beq"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup bge_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "bge";
    cp_asm_count : coverpoint ins.ins_str == "bge"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup bgeu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "bgeu";
    cp_asm_count : coverpoint ins.ins_str == "bgeu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup blt_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "blt";
    cp_asm_count : coverpoint ins.ins_str == "blt"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup bltu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "bltu";
    cp_asm_count : coverpoint ins.ins_str == "bltu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup bne_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "bne";
    cp_asm_count : coverpoint ins.ins_str == "bne"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_offset : coverpoint int'(ins.current.imm) - ins.get_pc()  iff (ins.trap == 0 )  {
        option.comment = "Branch Immediate Offset value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup jal_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "jal";
    cp_asm_count : coverpoint ins.ins_str == "jal"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rd_toggle_jal : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits. It has to be in multiples of 4. Therefore bit_0_1 and bit_1_1 are removed.";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }    cp_imm_ones_zeros_jal : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros. It has to be in multiples of 4. Therefore bit_0_1 and bit_1_1 are removed.";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup jalr_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "jalr";
    cp_asm_count : coverpoint ins.ins_str == "jalr"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rd_toggle_jal : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits. It has to be in multiples of 4. Therefore bit_0_1 and bit_1_1 are removed.";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup lb_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lb";
    cp_asm_count : coverpoint ins.ins_str == "lb"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rd_corners_lb : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111111111111111111111111111110000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111111111111111111111111111110000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000000000001111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000000000001111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111111111111111111111111111110101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000000000000000000000000000001010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000000000001011011};
        wildcard bins random1  = {64'b1111111111111111111111111111111111111111111111111111111111011011}; 
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup lbu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lbu";
    cp_asm_count : coverpoint ins.ins_str == "lbu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rd_corners_lbu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b0000000000000000000000000000000000000000000000000000000010000000};
        wildcard bins minp1    = {64'b0000000000000000000000000000000000000000000000000000000010000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000000000001111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000000000001111110};
        wildcard bins ones     = {64'b0000000000000000000000000000000000000000000000000000000011111111};
        wildcard bins onesm1   = {64'b0000000000000000000000000000000000000000000000000000000011111110};
        wildcard bins walkeodd = {64'b0000000000000000000000000000000000000000000000000000000010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000000000000000000000000000001010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000000000001011011};
        wildcard bins random1  = {64'b0000000000000000000000000000000000000000000000000000000011011011};  
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle_lbu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup ld_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "ld";
    cp_asm_count : coverpoint ins.ins_str == "ld"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
    cp_rd_boolean : coverpoint longint'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
endgroup

covergroup lh_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lh";
    cp_asm_count : coverpoint ins.ins_str == "lh"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
cp_rd_corners_lh : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111111111111111111111000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111111111111111111111000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b0000000000000000000000000000000000000000000000000101010101010101};
        wildcard bins walkeven = {64'b1111111111111111111111111111111111111111111111111010101010101010};
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000101101110111100};
        wildcard bins random1  = {64'b1111111111111111111111111111111111111111111111111101101110111100};
     }    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup lhu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lhu";
    cp_asm_count : coverpoint ins.ins_str == "lhu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
cp_rd_corners_lhu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0)  {
        option.comment = "RD Corners";
        wildcard bins zero     = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b0000000000000000000000000000000000000000000000001000000000000000};        // Zero Extended min half word
        wildcard bins minp1    = {64'b0000000000000000000000000000000000000000000000001000000000000001};        // Zero Extended minp1 half word
        wildcard bins max      = {64'b0000000000000000000000000000000000000000000000000111111111111111};        // Zero Extended max half word
        wildcard bins maxm1    = {64'b0000000000000000000000000000000000000000000000000111111111111110};        // Zero Extended maxm1 half word
        wildcard bins ones     = {64'b0000000000000000000000000000000000000000000000001111111111111111};        // Zero Extended ones half word
        wildcard bins onesm1   = {64'b0000000000000000000000000000000000000000000000001111111111111110};        // Zero Extended onesm1 half word
        wildcard bins walkeodd = {64'b0000000000000000000000000000000000000000000000000101010101010101};        // Zero Extended walkodd
        wildcard bins walkeven = {64'b0000000000000000000000000000000000000000000000001010101010101010};        // Zero Extended walkeven
        wildcard bins random0  = {64'b0000000000000000000000000000000000000000000000000101101110111100};        // Zero Extended random1
        wildcard bins random1  = {64'b0000000000000000000000000000000000000000000000001101101110111100};        // Zero Extended random1
     }    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle_lhu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup lui_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lui";
    cp_asm_count : coverpoint ins.ins_str == "lui"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
cp_rd_corners_lui : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0)  {
    option.comment = "RD Corners";
    wildcard bins zero   = {0};
    wildcard bins upper1 = {64'b1111111111111111111111111111111111111111111111111111000000000000};
    wildcard bins msb1   = {64'b1111111111111111111111111111111110000000000000000000000000000000};
    wildcard bins lsb1   = {64'b0000000000000000000000000000000000000000000000000001000000000000};
    wildcard bins random = {64'b0000000000000000000000000000000001001010111000100000000000000000};       
}
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm_zero : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate values";
        bins zero  = {0};
        bins nonzero  = default;
    }
endgroup

covergroup lw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lw";
    cp_asm_count : coverpoint ins.ins_str == "lw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
 cp_rd_corners_lw : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup lwu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "lwu";
    cp_asm_count : coverpoint ins.ins_str == "lwu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
 cp_rd_corners_lwu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b0000000000000000000000000000000010000000000000000000000000000000};
        wildcard bins minp1    = {64'b0000000000000000000000000000000010000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins onesm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins walkeodd = {64'b0000000000000000000000000000000010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b0000000000000000000000000000000011100011101011101000011011110111};
     }    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle_lwu : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_mem_hazard : coverpoint check_mem_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "Memory Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD};
    }
endgroup

covergroup or_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "or";
    cp_asm_count : coverpoint ins.ins_str == "or"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup ori_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "ori";
    cp_asm_count : coverpoint ins.ins_str == "ori"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup sb_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sb";
    cp_asm_count : coverpoint ins.ins_str == "sb"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup sd_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sd";
    cp_asm_count : coverpoint ins.ins_str == "sd"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup sh_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sh";
    cp_asm_count : coverpoint ins.ins_str == "sh"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup sll_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sll";
    cp_asm_count : coverpoint ins.ins_str == "sll"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup slli_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "slli";
    cp_asm_count : coverpoint ins.ins_str == "slli"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:63]};
    }
endgroup

covergroup slliw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "slliw";
    cp_asm_count : coverpoint ins.ins_str == "slliw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift_w : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift for W";
        bins shift[]  = {[0:31]};
    }
endgroup

covergroup sllw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sllw";
    cp_asm_count : coverpoint ins.ins_str == "sllw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup slt_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "slt";
    cp_asm_count : coverpoint ins.ins_str == "slt"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rd_boolean : coverpoint longint'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
endgroup

covergroup slti_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "slti";
    cp_asm_count : coverpoint ins.ins_str == "slti"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rd_boolean : coverpoint longint'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup sltiu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sltiu";
    cp_asm_count : coverpoint ins.ins_str == "sltiu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rd_boolean : coverpoint longint'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

covergroup sltu_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sltu";
    cp_asm_count : coverpoint ins.ins_str == "sltu"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rd_boolean : coverpoint longint'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Boolean Values";
        bins zero  = {0};
        bins one  = {1};
    }
endgroup

covergroup sra_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sra";
    cp_asm_count : coverpoint ins.ins_str == "sra"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup srai_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "srai";
    cp_asm_count : coverpoint ins.ins_str == "srai"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:63]};
    }
endgroup

covergroup sraiw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sraiw";
    cp_asm_count : coverpoint ins.ins_str == "sraiw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift_w : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift for W";
        bins shift[]  = {[0:31]};
    }
endgroup

covergroup sraw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sraw";
    cp_asm_count : coverpoint ins.ins_str == "sraw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup srl_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "srl";
    cp_asm_count : coverpoint ins.ins_str == "srl"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup srli_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "srli";
    cp_asm_count : coverpoint ins.ins_str == "srli"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift";
        bins shift[]  = {[0:63]};
    }
endgroup

covergroup srliw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "srliw";
    cp_asm_count : coverpoint ins.ins_str == "srliw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_shift_w : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate Shift for W";
        bins shift[]  = {[0:31]};
    }
endgroup

covergroup srlw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "srlw";
    cp_asm_count : coverpoint ins.ins_str == "srlw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup sub_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sub";
    cp_asm_count : coverpoint ins.ins_str == "sub"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup subw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "subw";
    cp_asm_count : coverpoint ins.ins_str == "subw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
   cp_rd_corners_32bit : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1111111111111111111111111111111110000000000000000000000000000000};
        wildcard bins minp1    = {64'b1111111111111111111111111111111110000000000000000000000000000001}; 
        wildcard bins max      = {64'b0000000000000000000000000000000001111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0000000000000000000000000000000001111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1111111111111111111111111111111110101010101010101010101010101010};
        wildcard bins walkeven = {64'b0000000000000000000000000000000001010101010101010101010101010101};
        wildcard bins random0  = {64'b0000000000000000000000000000000001100011101011101000011011110111};
        wildcard bins random1  = {64'b1111111111111111111111111111111111100011101011101000011011110111};
     }    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup sw_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "sw";
    cp_asm_count : coverpoint ins.ins_str == "sw"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rs1_nx0 : coverpoint ins.get_gpr_reg(ins.current.rs1) iff (ins.trap == 0) {
        option.comment = "RS1 register assignment (excluding x0)";

        bins x1 = {1};
        bins x2 = {2};
        bins x3 = {3};
        bins x4 = {4};
        bins x5 = {5};
        bins x6 = {6};
        bins x7 = {7};
        bins x8 = {8};
        bins x9 = {9};
        bins x10 = {10};
        bins x11 = {11};
        bins x12 = {12};
        bins x13 = {13};
        bins x14 = {14};
        bins x15 = {15};
        `ifndef COVER_BASE_E
        bins x16 = {16};
        bins x17 = {17};
        bins x18 = {18};
        bins x19 = {19};
        bins x20 = {20};
        bins x21 = {21};
        bins x22 = {22};
        bins x23 = {23};
        bins x24 = {24};
        bins x25 = {25};
        bins x26 = {26};
        bins x27 = {27};
        bins x28 = {28};
        bins x29 = {29};
        bins x30 = {30};
        bins x31 = {31};
        `endif    
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
endgroup

covergroup xor_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "xor";
    cp_asm_count : coverpoint ins.ins_str == "xor"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cp_rs2 : coverpoint ins.get_gpr_reg(ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RS2 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cmp_rd_rs2_eqval : coverpoint ins.current.rd_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS2 register values";
        bins rd_eqval_rs2  = {1};
        bins rd_neval_rs2  = {0};
    }
    cmp_rs1_rs2_eqval : coverpoint ins.current.rs1_val == ins.current.rs2_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register values";
        bins rs1_eqval_rs2  = {1};
        bins rs1_neval_rs2  = {0};
    }
    cp_gpr_hazard : coverpoint check_gpr_hazards(ins.hart, ins.issue)  iff (ins.trap == 0 )  {
        option.comment = "GPR Hazard";
        bins hazards[]  = {NO_HAZARD, RAW_HAZARD, WAR_HAZARD, WAW_HAZARD};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cp_rs2_corners : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cr_rs1_rs2_corners : cross cp_rs1_corners,cp_rs2_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 corners and RS2 corners";
    }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs2 : coverpoint ins.current.rd == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "RD and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rd_rs1_rs2 : coverpoint (ins.current.rd == ins.current.rs1) & (ins.current.rd == ins.current.rs2)  iff (ins.trap == 0 )  {
        option.comment = "RD, RS1, and RS2 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cmp_rs1_rs2 : coverpoint ins.current.rs1 == ins.current.rs2  iff (ins.trap == 0 )  {
        option.comment = "Compare RS1 and RS2 register assignment";
        bins x0  = {1} iff (ins.current.rs1 == "x0");
        bins x1  = {1} iff (ins.current.rs1 == "x1");
        bins x2  = {1} iff (ins.current.rs1 == "x2");
        bins x3  = {1} iff (ins.current.rs1 == "x3");
        bins x4  = {1} iff (ins.current.rs1 == "x4");
        bins x5  = {1} iff (ins.current.rs1 == "x5");
        bins x6  = {1} iff (ins.current.rs1 == "x6");
        bins x7  = {1} iff (ins.current.rs1 == "x7");
        bins x8  = {1} iff (ins.current.rs1 == "x8");
        bins x9  = {1} iff (ins.current.rs1 == "x9");
        bins x10  = {1} iff (ins.current.rs1 == "x10");
        bins x11  = {1} iff (ins.current.rs1 == "x11");
        bins x12  = {1} iff (ins.current.rs1 == "x12");
        bins x13  = {1} iff (ins.current.rs1 == "x13");
        bins x14  = {1} iff (ins.current.rs1 == "x14");
        bins x15  = {1} iff (ins.current.rs1 == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rs1 == "x16");
        bins x17  = {1} iff (ins.current.rs1 == "x17");
        bins x18  = {1} iff (ins.current.rs1 == "x18");
        bins x19  = {1} iff (ins.current.rs1 == "x19");
        bins x20  = {1} iff (ins.current.rs1 == "x20");
        bins x21  = {1} iff (ins.current.rs1 == "x21");
        bins x22  = {1} iff (ins.current.rs1 == "x22");
        bins x23  = {1} iff (ins.current.rs1 == "x23");
        bins x24  = {1} iff (ins.current.rs1 == "x24");
        bins x25  = {1} iff (ins.current.rs1 == "x25");
        bins x26  = {1} iff (ins.current.rs1 == "x26");
        bins x27  = {1} iff (ins.current.rs1 == "x27");
        bins x28  = {1} iff (ins.current.rs1 == "x28");
        bins x29  = {1} iff (ins.current.rs1 == "x29");
        bins x30  = {1} iff (ins.current.rs1 == "x30");
        bins x31  = {1} iff (ins.current.rs1 == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs2_sign : coverpoint int'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cr_rs1_rs2 : cross cp_rs1_sign,cp_rs2_sign  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and RS2 sign";
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs2_toggle : coverpoint unsigned'(ins.current.rs2_val)  iff (ins.trap == 0 )  {
        option.comment = "RS2 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
endgroup

covergroup xori_cg with function sample(ins_rv64i_t ins);
    option.per_instance = 1; 
    option.comment = "xori";
    cp_asm_count : coverpoint ins.ins_str == "xori"  iff (ins.trap == 0 )  {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint ins.get_gpr_reg(ins.current.rd)  iff (ins.trap == 0 )  {
        option.comment = "RD register assignment";
    }
    cp_rs1 : coverpoint ins.get_gpr_reg(ins.current.rs1)  iff (ins.trap == 0 )  {
        option.comment = "RS1 register assignment";
    }
    cmp_rd_rs1_eqval : coverpoint ins.current.rd_val == ins.current.rs1_val  iff (ins.trap == 0 )  {
        option.comment = "Compare RD and RS1 register values";
        bins rd_eqval_rs1  = {1};
        bins rd_neval_rs1  = {0};
    }
    cp_rd_corners : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
    }
    cp_rs1_corners : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Corners";
        wildcard bins zero  = {0};
        wildcard bins one      = {64'b0000000000000000000000000000000000000000000000000000000000000001};
        wildcard bins two      = {64'b0000000000000000000000000000000000000000000000000000000000000010};
        wildcard bins min      = {64'b1000000000000000000000000000000000000000000000000000000000000000};
        wildcard bins minp1    = {64'b1000000000000000000000000000000000000000000000000000000000000001}; 
        wildcard bins Wmax     = {64'b0000000000000000000000000000000011111111111111111111111111111111};
        wildcard bins Wmaxm1   = {64'b0000000000000000000000000000000011111111111111111111111111111110};
        wildcard bins Wmaxp1   = {64'b0000000000000000000000000000000100000000000000000000000000000000}; 
        wildcard bins Wmaxp2   = {64'b0000000000000000000000000000000100000000000000000000000000000001}; 
        wildcard bins max      = {64'b0111111111111111111111111111111111111111111111111111111111111111}; 
        wildcard bins maxm1    = {64'b0111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins ones     = {64'b1111111111111111111111111111111111111111111111111111111111111111};
        wildcard bins onesm1   = {64'b1111111111111111111111111111111111111111111111111111111111111110};
        wildcard bins walkeodd = {64'b1010101010101010101010101010101010101010101010101010101010101010};
        wildcard bins walkeven = {64'b0101010101010101010101010101010101010101010101010101010101010101};
        wildcard bins random   = {64'b0101101110111100100010000111011101100011101011101000011011110111};
     }
    cmp_rd_rs1 : coverpoint ins.current.rd == ins.current.rs1  iff (ins.trap == 0 )  {
        option.comment = "RD and RS1 register (assignment) WAR Hazard";
        bins x0  = {1} iff (ins.current.rd == "x0");
        bins x1  = {1} iff (ins.current.rd == "x1");
        bins x2  = {1} iff (ins.current.rd == "x2");
        bins x3  = {1} iff (ins.current.rd == "x3");
        bins x4  = {1} iff (ins.current.rd == "x4");
        bins x5  = {1} iff (ins.current.rd == "x5");
        bins x6  = {1} iff (ins.current.rd == "x6");
        bins x7  = {1} iff (ins.current.rd == "x7");
        bins x8  = {1} iff (ins.current.rd == "x8");
        bins x9  = {1} iff (ins.current.rd == "x9");
        bins x10  = {1} iff (ins.current.rd == "x10");
        bins x11  = {1} iff (ins.current.rd == "x11");
        bins x12  = {1} iff (ins.current.rd == "x12");
        bins x13  = {1} iff (ins.current.rd == "x13");
        bins x14  = {1} iff (ins.current.rd == "x14");
        bins x15  = {1} iff (ins.current.rd == "x15");
`ifndef COVER_BASE_E
        bins x16  = {1} iff (ins.current.rd == "x16");
        bins x17  = {1} iff (ins.current.rd == "x17");
        bins x18  = {1} iff (ins.current.rd == "x18");
        bins x19  = {1} iff (ins.current.rd == "x19");
        bins x20  = {1} iff (ins.current.rd == "x20");
        bins x21  = {1} iff (ins.current.rd == "x21");
        bins x22  = {1} iff (ins.current.rd == "x22");
        bins x23  = {1} iff (ins.current.rd == "x23");
        bins x24  = {1} iff (ins.current.rd == "x24");
        bins x25  = {1} iff (ins.current.rd == "x25");
        bins x26  = {1} iff (ins.current.rd == "x26");
        bins x27  = {1} iff (ins.current.rd == "x27");
        bins x28  = {1} iff (ins.current.rd == "x28");
        bins x29  = {1} iff (ins.current.rd == "x29");
        bins x30  = {1} iff (ins.current.rd == "x30");
        bins x31  = {1} iff (ins.current.rd == "x31");
`endif
    }
    cp_rd_sign : coverpoint int'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rs1_sign : coverpoint int'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 sign of value";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_imm_sign : coverpoint int'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value sign";
        bins neg  = {[$:-1]};
        bins pos  = {[1:$]};
    }
    cp_rd_toggle : coverpoint unsigned'(ins.current.rd_val)  iff (ins.trap == 0 )  {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_rs1_toggle : coverpoint unsigned'(ins.current.rs1_val)  iff (ins.trap == 0 )  {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0   = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0   = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0   = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0   = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0   = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0   = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0   = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0   = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0   = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0   = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_13_0  = {64'b??????????????????????????????????????????????????0?????????????};
        wildcard bins bit_14_0  = {64'b?????????????????????????????????????????????????0??????????????};
        wildcard bins bit_15_0  = {64'b????????????????????????????????????????????????0???????????????};
        wildcard bins bit_16_0  = {64'b???????????????????????????????????????????????0????????????????};
        wildcard bins bit_17_0  = {64'b??????????????????????????????????????????????0?????????????????};
        wildcard bins bit_18_0  = {64'b?????????????????????????????????????????????0??????????????????};
        wildcard bins bit_19_0  = {64'b????????????????????????????????????????????0???????????????????};
        wildcard bins bit_20_0  = {64'b???????????????????????????????????????????0????????????????????};
        wildcard bins bit_21_0  = {64'b??????????????????????????????????????????0?????????????????????};
        wildcard bins bit_22_0  = {64'b?????????????????????????????????????????0??????????????????????};
        wildcard bins bit_23_0  = {64'b????????????????????????????????????????0???????????????????????};
        wildcard bins bit_24_0  = {64'b???????????????????????????????????????0????????????????????????};
        wildcard bins bit_25_0  = {64'b??????????????????????????????????????0?????????????????????????};
        wildcard bins bit_26_0  = {64'b?????????????????????????????????????0??????????????????????????};
        wildcard bins bit_27_0  = {64'b????????????????????????????????????0???????????????????????????};
        wildcard bins bit_28_0  = {64'b???????????????????????????????????0????????????????????????????};
        wildcard bins bit_29_0  = {64'b??????????????????????????????????0?????????????????????????????};
        wildcard bins bit_30_0  = {64'b?????????????????????????????????0??????????????????????????????};
        wildcard bins bit_31_0  = {64'b????????????????????????????????0???????????????????????????????};
        wildcard bins bit_32_0  = {64'b???????????????????????????????0????????????????????????????????};
        wildcard bins bit_33_0  = {64'b??????????????????????????????0?????????????????????????????????};
        wildcard bins bit_34_0  = {64'b?????????????????????????????0??????????????????????????????????};
        wildcard bins bit_35_0  = {64'b????????????????????????????0???????????????????????????????????};
        wildcard bins bit_36_0  = {64'b???????????????????????????0????????????????????????????????????};
        wildcard bins bit_37_0  = {64'b??????????????????????????0?????????????????????????????????????};
        wildcard bins bit_38_0  = {64'b?????????????????????????0??????????????????????????????????????};
        wildcard bins bit_39_0  = {64'b????????????????????????0???????????????????????????????????????};
        wildcard bins bit_40_0  = {64'b???????????????????????0????????????????????????????????????????};
        wildcard bins bit_41_0  = {64'b??????????????????????0?????????????????????????????????????????};
        wildcard bins bit_42_0  = {64'b?????????????????????0??????????????????????????????????????????};
        wildcard bins bit_43_0  = {64'b????????????????????0???????????????????????????????????????????};
        wildcard bins bit_44_0  = {64'b???????????????????0????????????????????????????????????????????};
        wildcard bins bit_45_0  = {64'b??????????????????0?????????????????????????????????????????????};
        wildcard bins bit_46_0  = {64'b?????????????????0??????????????????????????????????????????????};
        wildcard bins bit_47_0  = {64'b????????????????0???????????????????????????????????????????????};
        wildcard bins bit_48_0  = {64'b???????????????0????????????????????????????????????????????????};
        wildcard bins bit_49_0  = {64'b??????????????0?????????????????????????????????????????????????};
        wildcard bins bit_50_0  = {64'b?????????????0??????????????????????????????????????????????????};
        wildcard bins bit_51_0  = {64'b????????????0???????????????????????????????????????????????????};
        wildcard bins bit_52_0  = {64'b???????????0????????????????????????????????????????????????????};
        wildcard bins bit_53_0  = {64'b??????????0?????????????????????????????????????????????????????};
        wildcard bins bit_54_0  = {64'b?????????0??????????????????????????????????????????????????????};
        wildcard bins bit_55_0  = {64'b????????0???????????????????????????????????????????????????????};
        wildcard bins bit_56_0  = {64'b???????0????????????????????????????????????????????????????????};
        wildcard bins bit_57_0  = {64'b??????0?????????????????????????????????????????????????????????};
        wildcard bins bit_58_0  = {64'b?????0??????????????????????????????????????????????????????????};
        wildcard bins bit_59_0  = {64'b????0???????????????????????????????????????????????????????????};
        wildcard bins bit_60_0  = {64'b???0????????????????????????????????????????????????????????????};
        wildcard bins bit_61_0  = {64'b??0?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_0  = {64'b?0??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_0  = {64'b0???????????????????????????????????????????????????????????????};
        wildcard bins bit_0_1   = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1   = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1   = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1   = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1   = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1   = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1   = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1   = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1   = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1   = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
        wildcard bins bit_13_1  = {64'b??????????????????????????????????????????????????1?????????????};
        wildcard bins bit_14_1  = {64'b?????????????????????????????????????????????????1??????????????};
        wildcard bins bit_15_1  = {64'b????????????????????????????????????????????????1???????????????};
        wildcard bins bit_16_1  = {64'b???????????????????????????????????????????????1????????????????};
        wildcard bins bit_17_1  = {64'b??????????????????????????????????????????????1?????????????????};
        wildcard bins bit_18_1  = {64'b?????????????????????????????????????????????1??????????????????};
        wildcard bins bit_19_1  = {64'b????????????????????????????????????????????1???????????????????};
        wildcard bins bit_20_1  = {64'b???????????????????????????????????????????1????????????????????};
        wildcard bins bit_21_1  = {64'b??????????????????????????????????????????1?????????????????????};
        wildcard bins bit_22_1  = {64'b?????????????????????????????????????????1??????????????????????};
        wildcard bins bit_23_1  = {64'b????????????????????????????????????????1???????????????????????};
        wildcard bins bit_24_1  = {64'b???????????????????????????????????????1????????????????????????};
        wildcard bins bit_25_1  = {64'b??????????????????????????????????????1?????????????????????????};
        wildcard bins bit_26_1  = {64'b?????????????????????????????????????1??????????????????????????};
        wildcard bins bit_27_1  = {64'b????????????????????????????????????1???????????????????????????};
        wildcard bins bit_28_1  = {64'b???????????????????????????????????1????????????????????????????};
        wildcard bins bit_29_1  = {64'b??????????????????????????????????1?????????????????????????????};
        wildcard bins bit_30_1  = {64'b?????????????????????????????????1??????????????????????????????};
        wildcard bins bit_31_1  = {64'b????????????????????????????????1???????????????????????????????};
        wildcard bins bit_32_1  = {64'b???????????????????????????????1????????????????????????????????};
        wildcard bins bit_33_1  = {64'b??????????????????????????????1?????????????????????????????????};
        wildcard bins bit_34_1  = {64'b?????????????????????????????1??????????????????????????????????};
        wildcard bins bit_35_1  = {64'b????????????????????????????1???????????????????????????????????};
        wildcard bins bit_36_1  = {64'b???????????????????????????1????????????????????????????????????};
        wildcard bins bit_37_1  = {64'b??????????????????????????1?????????????????????????????????????};
        wildcard bins bit_38_1  = {64'b?????????????????????????1??????????????????????????????????????};
        wildcard bins bit_39_1  = {64'b????????????????????????1???????????????????????????????????????};
        wildcard bins bit_40_1  = {64'b???????????????????????1????????????????????????????????????????};
        wildcard bins bit_41_1  = {64'b??????????????????????1?????????????????????????????????????????};
        wildcard bins bit_42_1  = {64'b?????????????????????1??????????????????????????????????????????};
        wildcard bins bit_43_1  = {64'b????????????????????1???????????????????????????????????????????};
        wildcard bins bit_44_1  = {64'b???????????????????1????????????????????????????????????????????};
        wildcard bins bit_45_1  = {64'b??????????????????1?????????????????????????????????????????????};
        wildcard bins bit_46_1  = {64'b?????????????????1??????????????????????????????????????????????};
        wildcard bins bit_47_1  = {64'b????????????????1???????????????????????????????????????????????};
        wildcard bins bit_48_1  = {64'b???????????????1????????????????????????????????????????????????};
        wildcard bins bit_49_1  = {64'b??????????????1?????????????????????????????????????????????????};
        wildcard bins bit_50_1  = {64'b?????????????1??????????????????????????????????????????????????};
        wildcard bins bit_51_1  = {64'b????????????1???????????????????????????????????????????????????};
        wildcard bins bit_52_1  = {64'b???????????1????????????????????????????????????????????????????};
        wildcard bins bit_53_1  = {64'b??????????1?????????????????????????????????????????????????????};
        wildcard bins bit_54_1  = {64'b?????????1??????????????????????????????????????????????????????};
        wildcard bins bit_55_1  = {64'b????????1???????????????????????????????????????????????????????};
        wildcard bins bit_56_1  = {64'b???????1????????????????????????????????????????????????????????};
        wildcard bins bit_57_1  = {64'b??????1?????????????????????????????????????????????????????????};
        wildcard bins bit_58_1  = {64'b?????1??????????????????????????????????????????????????????????};
        wildcard bins bit_59_1  = {64'b????1???????????????????????????????????????????????????????????};
        wildcard bins bit_60_1  = {64'b???1????????????????????????????????????????????????????????????};
        wildcard bins bit_61_1  = {64'b??1?????????????????????????????????????????????????????????????};
        wildcard bins bit_62_1  = {64'b?1??????????????????????????????????????????????????????????????};
        wildcard bins bit_63_1  = {64'b1???????????????????????????????????????????????????????????????};
    }
    cp_imm_ones_zeros : coverpoint unsigned'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Immediate value ones and zeros";
        wildcard bins bit_0_0  = {64'b???????????????????????????????????????????????????????????????0};
        wildcard bins bit_1_0  = {64'b??????????????????????????????????????????????????????????????0?};
        wildcard bins bit_2_0  = {64'b?????????????????????????????????????????????????????????????0??};
        wildcard bins bit_3_0  = {64'b????????????????????????????????????????????????????????????0???};
        wildcard bins bit_4_0  = {64'b???????????????????????????????????????????????????????????0????};
        wildcard bins bit_5_0  = {64'b??????????????????????????????????????????????????????????0?????};
        wildcard bins bit_6_0  = {64'b?????????????????????????????????????????????????????????0??????};
        wildcard bins bit_7_0  = {64'b????????????????????????????????????????????????????????0???????};
        wildcard bins bit_8_0  = {64'b???????????????????????????????????????????????????????0????????};
        wildcard bins bit_9_0  = {64'b??????????????????????????????????????????????????????0?????????};
        wildcard bins bit_10_0  = {64'b?????????????????????????????????????????????????????0??????????};
        wildcard bins bit_11_0  = {64'b????????????????????????????????????????????????????0???????????};
        wildcard bins bit_12_0  = {64'b???????????????????????????????????????????????????0????????????};
        wildcard bins bit_0_1  = {64'b???????????????????????????????????????????????????????????????1};
        wildcard bins bit_1_1  = {64'b??????????????????????????????????????????????????????????????1?};
        wildcard bins bit_2_1  = {64'b?????????????????????????????????????????????????????????????1??};
        wildcard bins bit_3_1  = {64'b????????????????????????????????????????????????????????????1???};
        wildcard bins bit_4_1  = {64'b???????????????????????????????????????????????????????????1????};
        wildcard bins bit_5_1  = {64'b??????????????????????????????????????????????????????????1?????};
        wildcard bins bit_6_1  = {64'b?????????????????????????????????????????????????????????1??????};
        wildcard bins bit_7_1  = {64'b????????????????????????????????????????????????????????1???????};
        wildcard bins bit_8_1  = {64'b???????????????????????????????????????????????????????1????????};
        wildcard bins bit_9_1  = {64'b??????????????????????????????????????????????????????1?????????};
        wildcard bins bit_10_1  = {64'b?????????????????????????????????????????????????????1??????????};
        wildcard bins bit_11_1  = {64'b????????????????????????????????????????????????????1???????????};
        wildcard bins bit_12_1  = {64'b???????????????????????????????????????????????????1????????????};
    }
    cp_imm12_corners : coverpoint signed'(ins.current.imm)  iff (ins.trap == 0 )  {
        option.comment = "Imm Corners";
        wildcard bins zero  = {0};
        wildcard bins one   = {1};
        wildcard bins two   = {2};
        wildcard bins hm1   = {1023};
        wildcard bins h   =   {1024};
        wildcard bins max   = {2047};
        wildcard bins min   = {-2048};
        wildcard bins minp1 = {-2047};
        wildcard bins onesm1 = {-2};
        wildcard bins ones  = {-1};
    }
    cr_rs1_imm_corners : cross cp_rs1_corners,cp_imm12_corners  iff (ins.trap == 0 )  {
        option.comment = "Cross coverage of RS1 sign and Imm corners";
    }
endgroup

function void rv64i_sample(int hart, int issue);
    ins_rv64i_t ins;

    case (traceDataQ[hart][issue][0].inst_name)
        "add"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            add_cg.sample(ins); 
        end
        "addi"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            addi_cg.sample(ins); 
        end
        "addiw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            addiw_cg.sample(ins); 
        end
        "addw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            addw_cg.sample(ins); 
        end
        "and"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            and_cg.sample(ins); 
        end
        "andi"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            andi_cg.sample(ins); 
        end
        "auipc"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            auipc_cg.sample(ins); 
        end
        "beq"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            beq_cg.sample(ins); 
        end
        "bge"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bge_cg.sample(ins); 
        end
        "bgeu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bgeu_cg.sample(ins); 
        end
        "blt"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            blt_cg.sample(ins); 
        end
        "bltu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bltu_cg.sample(ins); 
        end
        "bne"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs1(0);
            ins.add_rs2(1);
            ins.add_imm_addr(2);
            bne_cg.sample(ins); 
        end
        "jal"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm_addr(1);
            jal_cg.sample(ins); 
        end
        "jalr"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            if (ins.ops[2].key) begin           // To handle the form (instr rd, imm(rs1))
                ins.add_imm_addr(1);
                ins.add_rs1(2);
            end else if (ins.ops[1].key) begin  // To handle the form (instr rd, rs1)
                ins.add_rs1(1);
            end else begin                      // To handle compressed form (instr rs1)
                ins.add_rd_1();
                ins.add_rs1(0);
            end
            jalr_cg.sample(ins); 
        end
        "lb"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lb_cg.sample(ins); 
        end
        "lbu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lbu_cg.sample(ins); 
        end
        "ld"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            ld_cg.sample(ins); 
        end
        "lh"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lh_cg.sample(ins); 
        end
        "lhu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lhu_cg.sample(ins); 
        end
        "lui"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            lui_cg.sample(ins); 
        end
        "lw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lw_cg.sample(ins); 
        end
        "lwu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_LOAD;
            ins.add_mem_address();
            lwu_cg.sample(ins); 
        end
        "or"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            or_cg.sample(ins); 
        end
        "ori"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            ori_cg.sample(ins); 
        end
        "sb"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sb_cg.sample(ins); 
        end
        "sd"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sd_cg.sample(ins); 
        end
        "sh"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sh_cg.sample(ins); 
        end
        "sll"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sll_cg.sample(ins); 
        end
        "slli"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            slli_cg.sample(ins); 
        end
        "slliw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            slliw_cg.sample(ins); 
        end
        "sllw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sllw_cg.sample(ins); 
        end
        "slt"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            slt_cg.sample(ins); 
        end
        "slti"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            slti_cg.sample(ins); 
        end
        "sltiu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            sltiu_cg.sample(ins); 
        end
        "sltu"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sltu_cg.sample(ins); 
        end
        "sra"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sra_cg.sample(ins); 
        end
        "srai"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            srai_cg.sample(ins); 
        end
        "sraiw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            sraiw_cg.sample(ins); 
        end
        "sraw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sraw_cg.sample(ins); 
        end
        "srl"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            srl_cg.sample(ins); 
        end
        "srli"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            srli_cg.sample(ins); 
        end
        "srliw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            srliw_cg.sample(ins); 
        end
        "srlw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            srlw_cg.sample(ins); 
        end
        "sub"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            sub_cg.sample(ins); 
        end
        "subw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            subw_cg.sample(ins); 
        end
        "sw"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rs2(0);
            ins.add_imm(1);
            ins.add_rs1(2);
            ins.current.inst_category = INST_CAT_STORE;
            ins.add_mem_address();
            sw_cg.sample(ins); 
        end
        "xor"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_rs2(2);
            xor_cg.sample(ins); 
        end
        "xori"     : begin 
            ins = new(hart, issue, traceDataQ); 
            ins.add_rd(0);
            ins.add_rs1(1);
            ins.add_imm(2);
            xori_cg.sample(ins); 
        end
    endcase
endfunction
