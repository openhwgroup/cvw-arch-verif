///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    ZicsrS_scause_cg = new();      ZicsrS_scause_cg.set_inst_name("obj_scause");
    ZicsrS_sstatus_cg = new();     ZicsrS_sstatus_cg.set_inst_name("obj_sstatus");
    ZicsrS_sprivinst_cg = new();   ZicsrS_sprivinst_cg.set_inst_name("obj_sprivinst");
