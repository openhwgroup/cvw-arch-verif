///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////
    Svinval_sfence_inval_ir_cg = new(); Svinval_sfence_inval_ir_cg.set_inst_name("obj_Svinval_sfence_inval_ir");
    Svinval_sfence_w_inval_cg = new(); Svinval_sfence_w_inval_cg.set_inst_name("obj_Svinval_sfence_w_inval");
    Svinval_sinval_vma_cg = new(); Svinval_sinval_vma_cg.set_inst_name("obj_Svinval_sinval_vma");
