///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_ZICSRF
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_zicsrf_t;

covergroup fcsr_cg with function sample(ins_zicsrf_t ins);
    option.per_instance = 1; 
    option.comment = "ZicsrF fcsr";

    // building blocks for the main coverpoints

    csrrw_fcsr: coverpoint ins.current.insn {
        wildcard bins csrrw_fcsr = {32'b000000000011_?????_001_?????_1110011}; 
    }
    fcsr_frm_corners: coverpoint ins.current.rs1_val[7:5] {

    }
    fflags_corners: coverpoint ins.current.rs1_val[4:0] {

    }
    fcsr_reserved_walking: coverpoint ins.current.rs1_val[(XLEN-1):8]{
        `ifdef XLEN64
        bins b_8  = {56'b00000000000000000000000000000000000000000000000000000001};
        bins b_9  = {56'b00000000000000000000000000000000000000000000000000000010};
        bins b_10 = {56'b00000000000000000000000000000000000000000000000000000100};
        bins b_11 = {56'b00000000000000000000000000000000000000000000000000001000};
        bins b_12 = {56'b00000000000000000000000000000000000000000000000000010000};
        bins b_13 = {56'b00000000000000000000000000000000000000000000000000100000};
        bins b_14 = {56'b00000000000000000000000000000000000000000000000001000000};
        bins b_15 = {56'b00000000000000000000000000000000000000000000000010000000};
        bins b_16 = {56'b00000000000000000000000000000000000000000000000100000000};
        bins b_17 = {56'b00000000000000000000000000000000000000000000001000000000};
        bins b_18 = {56'b00000000000000000000000000000000000000000000010000000000};
        bins b_19 = {56'b00000000000000000000000000000000000000000000100000000000};
        bins b_20 = {56'b00000000000000000000000000000000000000000001000000000000};
        bins b_21 = {56'b00000000000000000000000000000000000000000010000000000000};
        bins b_22 = {56'b00000000000000000000000000000000000000000100000000000000};
        bins b_23 = {56'b00000000000000000000000000000000000000001000000000000000};
        bins b_24 = {56'b00000000000000000000000000000000000000010000000000000000};
        bins b_25 = {56'b00000000000000000000000000000000000000100000000000000000};
        bins b_26 = {56'b00000000000000000000000000000000000001000000000000000000};
        bins b_27 = {56'b00000000000000000000000000000000000010000000000000000000};
        bins b_28 = {56'b00000000000000000000000000000000000100000000000000000000};
        bins b_29 = {56'b00000000000000000000000000000000001000000000000000000000};
        bins b_30 = {56'b00000000000000000000000000000000010000000000000000000000};
        bins b_31 = {56'b00000000000000000000000000000000100000000000000000000000};
        bins b_32 = {56'b00000000000000000000000000000001000000000000000000000000};
        bins b_33 = {56'b00000000000000000000000000000010000000000000000000000000};
        bins b_34 = {56'b00000000000000000000000000000100000000000000000000000000};
        bins b_35 = {56'b00000000000000000000000000001000000000000000000000000000};
        bins b_36 = {56'b00000000000000000000000000010000000000000000000000000000};
        bins b_37 = {56'b00000000000000000000000000100000000000000000000000000000};
        bins b_38 = {56'b00000000000000000000000001000000000000000000000000000000};
        bins b_39 = {56'b00000000000000000000000010000000000000000000000000000000};
        bins b_40 = {56'b00000000000000000000000100000000000000000000000000000000};
        bins b_41 = {56'b00000000000000000000001000000000000000000000000000000000};
        bins b_42 = {56'b00000000000000000000010000000000000000000000000000000000};
        bins b_43 = {56'b00000000000000000000100000000000000000000000000000000000};
        bins b_44 = {56'b00000000000000000001000000000000000000000000000000000000};
        bins b_45 = {56'b00000000000000000010000000000000000000000000000000000000};
        bins b_46 = {56'b00000000000000000100000000000000000000000000000000000000};
        bins b_47 = {56'b00000000000000001000000000000000000000000000000000000000};
        bins b_48 = {56'b00000000000000010000000000000000000000000000000000000000};
        bins b_49 = {56'b00000000000000100000000000000000000000000000000000000000};
        bins b_50 = {56'b00000000000001000000000000000000000000000000000000000000};
        bins b_51 = {56'b00000000000010000000000000000000000000000000000000000000};
        bins b_52 = {56'b00000000000100000000000000000000000000000000000000000000};
        bins b_53 = {56'b00000000001000000000000000000000000000000000000000000000};
        bins b_54 = {56'b00000000010000000000000000000000000000000000000000000000};
        bins b_55 = {56'b00000000100000000000000000000000000000000000000000000000};
        bins b_56 = {56'b00000001000000000000000000000000000000000000000000000000};
        bins b_57 = {56'b00000010000000000000000000000000000000000000000000000000};
        bins b_58 = {56'b00000100000000000000000000000000000000000000000000000000};
        bins b_59 = {56'b00001000000000000000000000000000000000000000000000000000};
        bins b_60 = {56'b00010000000000000000000000000000000000000000000000000000};
        bins b_61 = {56'b00100000000000000000000000000000000000000000000000000000};
        bins b_62 = {56'b01000000000000000000000000000000000000000000000000000000};
        bins b_63 = {56'b10000000000000000000000000000000000000000000000000000000};
        `else
        bins b_8  = {24'b000000000000000000000001};
        bins b_9  = {24'b000000000000000000000010};
        bins b_10 = {24'b000000000000000000000100};
        bins b_11 = {24'b000000000000000000001000};
        bins b_12 = {24'b000000000000000000010000};
        bins b_13 = {24'b000000000000000000100000};
        bins b_14 = {24'b000000000000000001000000};
        bins b_15 = {24'b000000000000000010000000};
        bins b_16 = {24'b000000000000000100000000};
        bins b_17 = {24'b000000000000001000000000};
        bins b_18 = {24'b000000000000010000000000};
        bins b_19 = {24'b000000000000100000000000};
        bins b_20 = {24'b000000000001000000000000};
        bins b_21 = {24'b000000000010000000000000};
        bins b_22 = {24'b000000000100000000000000};
        bins b_23 = {24'b000000001000000000000000};
        bins b_24 = {24'b000000010000000000000000};
        bins b_25 = {24'b000000100000000000000000};
        bins b_26 = {24'b000001000000000000000000};
        bins b_27 = {24'b000010000000000000000000};
        bins b_28 = {24'b000100000000000000000000};
        bins b_29 = {24'b001000000000000000000000};
        bins b_30 = {24'b010000000000000000000000};
        bins b_31 = {24'b100000000000000000000000};
        `endif
    }
    mstatus_FS: coverpoint ins.current.csr[12'h300][14:13] {

    }
    
    // main coverpoints
    cp_fcsr_frm_write:    cross csrrw_fcsr, fcsr_frm_corners,      mstatus_FS;
    cp_fcsr_fflags_write: cross csrrw_fcsr, fflags_corners,        mstatus_FS;
    cp_fcsr_reserved:     cross csrrw_fcsr, fcsr_reserved_walking, mstatus_FS; 
endgroup

covergroup frm_cg with function sample(ins_zicsrf_t ins);
    option.per_instance = 1; 
    option.comment = "ZicsrF frm csr";

    // building blocks for main coverpoints
    csrrw_frm: coverpoint ins.current.insn {
    wildcard bins csrrw_frm = {32'b000000000010_?????_001_?????_1110011}; 
    }
    frm_corners: coverpoint ins.current.rs1_val[2:0] {

    }
    frm_reserved_walking: coverpoint ins.current.rs1_val[(XLEN-1):3] {
        `ifdef XLEN64
        bins b_3  = {61'b0000000000000000000000000000000000000000000000000000000000001};
        bins b_4  = {61'b0000000000000000000000000000000000000000000000000000000000010};
        bins b_5  = {61'b0000000000000000000000000000000000000000000000000000000000100};
        bins b_6  = {61'b0000000000000000000000000000000000000000000000000000000001000};
        bins b_7  = {61'b0000000000000000000000000000000000000000000000000000000010000};
        bins b_8  = {61'b0000000000000000000000000000000000000000000000000000000100000};
        bins b_9  = {61'b0000000000000000000000000000000000000000000000000000001000000};
        bins b_10 = {61'b0000000000000000000000000000000000000000000000000000010000000};
        bins b_11 = {61'b0000000000000000000000000000000000000000000000000000100000000};
        bins b_12 = {61'b0000000000000000000000000000000000000000000000000001000000000};
        bins b_13 = {61'b0000000000000000000000000000000000000000000000000010000000000};
        bins b_14 = {61'b0000000000000000000000000000000000000000000000000100000000000};
        bins b_15 = {61'b0000000000000000000000000000000000000000000000001000000000000};
        bins b_16 = {61'b0000000000000000000000000000000000000000000000010000000000000};
        bins b_17 = {61'b0000000000000000000000000000000000000000000000100000000000000};
        bins b_18 = {61'b0000000000000000000000000000000000000000000001000000000000000};
        bins b_19 = {61'b0000000000000000000000000000000000000000000010000000000000000};
        bins b_20 = {61'b0000000000000000000000000000000000000000000100000000000000000};
        bins b_21 = {61'b0000000000000000000000000000000000000000001000000000000000000};
        bins b_22 = {61'b0000000000000000000000000000000000000000010000000000000000000};
        bins b_23 = {61'b0000000000000000000000000000000000000000100000000000000000000};
        bins b_24 = {61'b0000000000000000000000000000000000000001000000000000000000000};
        bins b_25 = {61'b0000000000000000000000000000000000000010000000000000000000000};
        bins b_26 = {61'b0000000000000000000000000000000000000100000000000000000000000};
        bins b_27 = {61'b0000000000000000000000000000000000001000000000000000000000000};
        bins b_28 = {61'b0000000000000000000000000000000000010000000000000000000000000};
        bins b_29 = {61'b0000000000000000000000000000000000100000000000000000000000000};
        bins b_30 = {61'b0000000000000000000000000000000001000000000000000000000000000};
        bins b_31 = {61'b0000000000000000000000000000000010000000000000000000000000000};
        bins b_32 = {61'b0000000000000000000000000000000100000000000000000000000000000};
        bins b_33 = {61'b0000000000000000000000000000001000000000000000000000000000000};
        bins b_34 = {61'b0000000000000000000000000000010000000000000000000000000000000};
        bins b_35 = {61'b0000000000000000000000000000100000000000000000000000000000000};
        bins b_36 = {61'b0000000000000000000000000001000000000000000000000000000000000};
        bins b_37 = {61'b0000000000000000000000000010000000000000000000000000000000000};
        bins b_38 = {61'b0000000000000000000000000100000000000000000000000000000000000};
        bins b_39 = {61'b0000000000000000000000001000000000000000000000000000000000000};
        bins b_40 = {61'b0000000000000000000000010000000000000000000000000000000000000};
        bins b_41 = {61'b0000000000000000000000100000000000000000000000000000000000000};
        bins b_42 = {61'b0000000000000000000001000000000000000000000000000000000000000};
        bins b_43 = {61'b0000000000000000000010000000000000000000000000000000000000000};
        bins b_44 = {61'b0000000000000000000100000000000000000000000000000000000000000};
        bins b_45 = {61'b0000000000000000001000000000000000000000000000000000000000000};
        bins b_46 = {61'b0000000000000000010000000000000000000000000000000000000000000};
        bins b_47 = {61'b0000000000000000100000000000000000000000000000000000000000000};
        bins b_48 = {61'b0000000000000001000000000000000000000000000000000000000000000};
        bins b_49 = {61'b0000000000000010000000000000000000000000000000000000000000000};
        bins b_50 = {61'b0000000000000100000000000000000000000000000000000000000000000};
        bins b_51 = {61'b0000000000001000000000000000000000000000000000000000000000000};
        bins b_52 = {61'b0000000000010000000000000000000000000000000000000000000000000};
        bins b_53 = {61'b0000000000100000000000000000000000000000000000000000000000000};
        bins b_54 = {61'b0000000001000000000000000000000000000000000000000000000000000};
        bins b_55 = {61'b0000000010000000000000000000000000000000000000000000000000000};
        bins b_56 = {61'b0000000100000000000000000000000000000000000000000000000000000};
        bins b_57 = {61'b0000001000000000000000000000000000000000000000000000000000000};
        bins b_58 = {61'b0000010000000000000000000000000000000000000000000000000000000};
        bins b_59 = {61'b0000100000000000000000000000000000000000000000000000000000000};
        bins b_60 = {61'b0001000000000000000000000000000000000000000000000000000000000};
        bins b_61 = {61'b0010000000000000000000000000000000000000000000000000000000000};
        bins b_62 = {61'b0100000000000000000000000000000000000000000000000000000000000};
        bins b_63 = {61'b1000000000000000000000000000000000000000000000000000000000000};
        `else 
        bins b_3  = {29'b00000000000000000000000000001};
        bins b_4  = {29'b00000000000000000000000000010};
        bins b_5  = {29'b00000000000000000000000000100};
        bins b_6  = {29'b00000000000000000000000001000};
        bins b_7  = {29'b00000000000000000000000010000};
        bins b_8  = {29'b00000000000000000000000100000};
        bins b_9  = {29'b00000000000000000000001000000};
        bins b_10 = {29'b00000000000000000000010000000};
        bins b_11 = {29'b00000000000000000000100000000};
        bins b_12 = {29'b00000000000000000001000000000};
        bins b_13 = {29'b00000000000000000010000000000};
        bins b_14 = {29'b00000000000000000100000000000};
        bins b_15 = {29'b00000000000000001000000000000};
        bins b_16 = {29'b00000000000000010000000000000};
        bins b_17 = {29'b00000000000000100000000000000};
        bins b_18 = {29'b00000000000001000000000000000};
        bins b_19 = {29'b00000000000010000000000000000};
        bins b_20 = {29'b00000000000100000000000000000};
        bins b_21 = {29'b00000000001000000000000000000};
        bins b_22 = {29'b00000000010000000000000000000};
        bins b_23 = {29'b00000000100000000000000000000};
        bins b_24 = {29'b00000001000000000000000000000};
        bins b_25 = {29'b00000010000000000000000000000};
        bins b_26 = {29'b00000100000000000000000000000};
        bins b_27 = {29'b00001000000000000000000000000};
        bins b_28 = {29'b00010000000000000000000000000};
        bins b_29 = {29'b00100000000000000000000000000};
        bins b_30 = {29'b01000000000000000000000000000};
        bins b_31 = {29'b10000000000000000000000000000};
        `endif
    }
    mstatus_FS: coverpoint ins.current.csr[12'h300][14:13] {

    }
    // main coverpoints
    cp_frm_write:          cross csrrw_frm, frm_corners,          mstatus_FS;
    cp_frm_write_reserved: cross csrrw_frm, frm_reserved_walking, mstatus_FS;
endgroup

covergroup fflags_cg with function sample(ins_zicsrf_t ins);
    option.per_instance = 1; 
    option.comment = "ZicsrF fflags csr";

    // building blocks for main coverpoints
    csrrw_fflags: coverpoint ins.current.insn {
    wildcard bins csrrw_fflags = {32'b000000000001_?????_001_?????_1110011}; 
    }
    fflags_corners: coverpoint ins.current.rs1_val[4:0] {

    }
    fflags_reserved_walking: coverpoint ins.current.rs1_val[(XLEN-1):5] {
        `ifdef XLEN64
        bins b_5  = {59'b00000000000000000000000000000000000000000000000000000000001};
        bins b_6  = {59'b00000000000000000000000000000000000000000000000000000000010};
        bins b_7  = {59'b00000000000000000000000000000000000000000000000000000000100};
        bins b_8  = {59'b00000000000000000000000000000000000000000000000000000001000};
        bins b_9  = {59'b00000000000000000000000000000000000000000000000000000010000};
        bins b_10 = {59'b00000000000000000000000000000000000000000000000000000100000};
        bins b_11 = {59'b00000000000000000000000000000000000000000000000000001000000};
        bins b_12 = {59'b00000000000000000000000000000000000000000000000000010000000};
        bins b_13 = {59'b00000000000000000000000000000000000000000000000000100000000};
        bins b_14 = {59'b00000000000000000000000000000000000000000000000001000000000};
        bins b_15 = {59'b00000000000000000000000000000000000000000000000010000000000};
        bins b_16 = {59'b00000000000000000000000000000000000000000000000100000000000};
        bins b_17 = {59'b00000000000000000000000000000000000000000000001000000000000};
        bins b_18 = {59'b00000000000000000000000000000000000000000000010000000000000};
        bins b_19 = {59'b00000000000000000000000000000000000000000000100000000000000};
        bins b_20 = {59'b00000000000000000000000000000000000000000001000000000000000};
        bins b_21 = {59'b00000000000000000000000000000000000000000010000000000000000};
        bins b_22 = {59'b00000000000000000000000000000000000000000100000000000000000};
        bins b_23 = {59'b00000000000000000000000000000000000000001000000000000000000};
        bins b_24 = {59'b00000000000000000000000000000000000000010000000000000000000};
        bins b_25 = {59'b00000000000000000000000000000000000000100000000000000000000};
        bins b_26 = {59'b00000000000000000000000000000000000001000000000000000000000};
        bins b_27 = {59'b00000000000000000000000000000000000010000000000000000000000};
        bins b_28 = {59'b00000000000000000000000000000000000100000000000000000000000};
        bins b_29 = {59'b00000000000000000000000000000000001000000000000000000000000};
        bins b_30 = {59'b00000000000000000000000000000000010000000000000000000000000};
        bins b_31 = {59'b00000000000000000000000000000000100000000000000000000000000};
        bins b_32 = {59'b00000000000000000000000000000001000000000000000000000000000};
        bins b_33 = {59'b00000000000000000000000000000010000000000000000000000000000};
        bins b_34 = {59'b00000000000000000000000000000100000000000000000000000000000};
        bins b_35 = {59'b00000000000000000000000000001000000000000000000000000000000};
        bins b_36 = {59'b00000000000000000000000000010000000000000000000000000000000};
        bins b_37 = {59'b00000000000000000000000000100000000000000000000000000000000};
        bins b_38 = {59'b00000000000000000000000001000000000000000000000000000000000};
        bins b_39 = {59'b00000000000000000000000010000000000000000000000000000000000};
        bins b_40 = {59'b00000000000000000000000100000000000000000000000000000000000};
        bins b_41 = {59'b00000000000000000000001000000000000000000000000000000000000};
        bins b_42 = {59'b00000000000000000000010000000000000000000000000000000000000};
        bins b_43 = {59'b00000000000000000000100000000000000000000000000000000000000};
        bins b_44 = {59'b00000000000000000001000000000000000000000000000000000000000};
        bins b_45 = {59'b00000000000000000010000000000000000000000000000000000000000};
        bins b_46 = {59'b00000000000000000100000000000000000000000000000000000000000};
        bins b_47 = {59'b00000000000000001000000000000000000000000000000000000000000};
        bins b_48 = {59'b00000000000000010000000000000000000000000000000000000000000};
        bins b_49 = {59'b00000000000000100000000000000000000000000000000000000000000};
        bins b_50 = {59'b00000000000001000000000000000000000000000000000000000000000};
        bins b_51 = {59'b00000000000010000000000000000000000000000000000000000000000};
        bins b_52 = {59'b00000000000100000000000000000000000000000000000000000000000};
        bins b_53 = {59'b00000000001000000000000000000000000000000000000000000000000};
        bins b_54 = {59'b00000000010000000000000000000000000000000000000000000000000};
        bins b_55 = {59'b00000000100000000000000000000000000000000000000000000000000};
        bins b_56 = {59'b00000001000000000000000000000000000000000000000000000000000};
        bins b_57 = {59'b00000010000000000000000000000000000000000000000000000000000};
        bins b_58 = {59'b00000100000000000000000000000000000000000000000000000000000};
        bins b_59 = {59'b00001000000000000000000000000000000000000000000000000000000};
        bins b_60 = {59'b00010000000000000000000000000000000000000000000000000000000};
        bins b_61 = {59'b00100000000000000000000000000000000000000000000000000000000};
        bins b_62 = {59'b01000000000000000000000000000000000000000000000000000000000};
        bins b_63 = {59'b10000000000000000000000000000000000000000000000000000000000};
        `else
        bins b_5  = {27'b000000000000000000000000001};
        bins b_6  = {27'b000000000000000000000000010};
        bins b_7  = {27'b000000000000000000000000100};
        bins b_8  = {27'b000000000000000000000001000};
        bins b_9  = {27'b000000000000000000000010000};
        bins b_10 = {27'b000000000000000000000100000};
        bins b_11 = {27'b000000000000000000001000000};
        bins b_12 = {27'b000000000000000000010000000};
        bins b_13 = {27'b000000000000000000100000000};
        bins b_14 = {27'b000000000000000001000000000};
        bins b_15 = {27'b000000000000000010000000000};
        bins b_16 = {27'b000000000000000100000000000};
        bins b_17 = {27'b000000000000001000000000000};
        bins b_18 = {27'b000000000000010000000000000};
        bins b_19 = {27'b000000000000100000000000000};
        bins b_20 = {27'b000000000001000000000000000};
        bins b_21 = {27'b000000000010000000000000000};
        bins b_22 = {27'b000000000100000000000000000};
        bins b_23 = {27'b000000001000000000000000000};
        bins b_24 = {27'b000000010000000000000000000};
        bins b_25 = {27'b000000100000000000000000000};
        bins b_26 = {27'b000001000000000000000000000};
        bins b_27 = {27'b000010000000000000000000000};
        bins b_28 = {27'b000100000000000000000000000};
        bins b_29 = {27'b001000000000000000000000000};
        bins b_30 = {27'b010000000000000000000000000};
        bins b_31 = {27'b100000000000000000000000000};
        `endif
    }
    fflags_toggle: coverpoint ins.current.csr[12'h003][4:0] {
        wildcard bins NX = (5'b????0 => 5'b????1);
        wildcard bins UF = (5'b???0? => 5'b???1?);
        wildcard bins OF = (5'b??0?? => 5'b??1??);
        wildcard bins DZ = (5'b?0??? => 5'b?1???);
        wildcard bins NV = (5'b0???? => 5'b1????);
    }
    mstatus_FS: coverpoint ins.current.csr[12'h300][14:13] {

    }
    mstatus_FS_n0: coverpoint ins.current.csr[12'h300][14:13] {
        bins not_zero = {!3'b000};
    }
    // main coverpoints
    cp_fflags_write:          cross csrrw_fflags, fflags_corners,          mstatus_FS;
    cp_fflags_write_reserved: cross csrrw_fflags, fflags_reserved_walking, mstatus_FS;
    cp_fflags_set_m:          cross fflags_toggle, mstatus_FS_n0;
endgroup

function void zicsrf_sample(int hart, int issue);
    ins_zicsrf_t ins;

    ins = new(hart, issue, traceDataQ); 
    ins.add_rd(0);
    ins.add_rs1(2);
    ins.add_csr(1);
    
    fcsr_cg.sample(ins);
    frm_cg.sample(ins);
    fflags_cg.sample(ins);
    
endfunction
