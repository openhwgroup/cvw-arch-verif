///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups
// 
// Written: David_Harris@hmc.edu 26 November 2024
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may not use this file 
// except in compliance with the License, or, at your option, the Apache License version 2.0. You 
// may obtain a copy of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work distributed under the 
// License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, 
// either express or implied. See the License for the specific language governing permissions 
// and limitations under the License.
////////////////////////////////////////////////////////////////////////////////////////////////

`define COVER_EXCEPTIONSINSTR
typedef RISCV_instruction #(ILEN, XLEN, FLEN, VLEN, NHART, RETIRE) ins_exceptionsinstr_t;

covergroup exceptionsInstr_cg with function sample(ins_exceptionsinstr_t ins);
    option.per_instance = 0; 
    
    cp_legalI : coverpoint ins.current.insn iff (ins.trap == 0 )  {
        wildcard bins lb = {32'b????????????_?????_000_?????_0000011};
        wildcard bins lh = {32'b????????????_?????_001_?????_0000011};
    }
    cp_illegal : coverpoint ins.current.insn iff (ins.trap == 1) { // should trap
    	wildcard bins op2  = {32'b?????????????????????????_0001011}; // unused ops
    	wildcard bins op7  = {32'b?????????????????????????_0011111}; // unused ops
    	wildcard bins op10 = {32'b?????????????????????????_0101011}; // unused ops
    	wildcard bins op15 = {32'b?????????????????????????_0111111}; // unused ops
    	wildcard bins op21 = {32'b?????????????????????????_1010111}; // unused ops
    	wildcard bins op22 = {32'b?????????????????????????_1011011}; // unused ops
    	wildcard bins op23 = {32'b?????????????????????????_1011111}; // unused ops
    	wildcard bins op26 = {32'b?????????????????????????_1101011}; // unused ops
    	wildcard bins op29 = {32'b?????????????????????????_1110111}; // unused ops
    	wildcard bins op30 = {32'b?????????????????????????_1111011}; // unused ops
    	wildcard bins op31 = {32'b?????????????????????????_1111111}; // unused ops
        // load instructions with illegal funct3
    	wildcard bins illegal_load = {32'b????????????_?????_111_00000_0000011}; // load with funct3 = 7
        `ifdef XLEN32
    	    wildcard bins illegal_ld =  {32'b????????????_?????_011_?????_0000011}; // ld
            wildcard bins illegal_lwu = {32'b????????????_?????_110_?????_0000011}; // lwu
        `endif
        // floating-point load instructions with illegal funct3
    	wildcard bins illegal_fload0 = {32'b????????????_?????_000_?????_0000111}; // fp load with funct3 = 0
    	wildcard bins illegal_fload0 = {32'b????????????_?????_101_?????_0000111}; // fp load with funct3 = 5
    	wildcard bins illegal_fload0 = {32'b????????????_?????_110_?????_0000111}; // fp load with funct3 = 6
    	wildcard bins illegal_fload0 = {32'b????????????_?????_111_?????_0000111}; // fp load with funct3 = 7
        // fence/cbo instructions with illegal funct3
    	wildcard bins illegal_fence3 = {32'b????????????_?????_011_?????_0001111}; // fence/cbo with funct3 = 3
        
    }

endgroup

function void exceptionsinstr_sample(int hart, int issue);
    ins_exceptionsinstr_t ins;

    ins = new(hart, issue, traceDataQ); 

//    $display("Instruction is: PC %h: %h = %s (rd = %h rs1 = %h rs2 = %h) trap = %b mode = %b (old mode %b) mstatus %h (old mstatus %h).  Retired: %d",ins.current.pc_rdata, ins.current.insn, ins.current.disass, ins.current.rd_val, ins.current.rs1_val, ins.current.rs2_val, ins.current.trap, ins.current.mode, ins.prev.mode, ins.current.csr[12'h300], ins.prev.csr[12'h300], ins.current.csr[12'hB02]);
//    $display("Instruction is: %b %b %s", ins.current.insn[14:12], ins.current.insn[6:0], ins.current.disass);
    
    exceptionsInstr_cg.sample(ins);
    
endfunction
