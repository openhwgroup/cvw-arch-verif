///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    aaes64es_cg = new(); aaes64es_cg.set_inst_name("obj_aaes64es");
    aes64esmi_cg = new(); aes64esmi_cg.set_inst_name("obj_aes64esmi");
    aes64ks1i_cg = new(); aes64ks1i_cg.set_inst_name("obj_aes64ks1i");
    aes64ks2_cg = new(); aes64ks2_cg.set_inst_name("obj_aes64ks2");
