///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    clmul_cg = new(); clmul_cg.set_inst_name("obj_clmul");
    clmulh_cg = new(); clmulh_cg.set_inst_name("obj_clmulh");
    clmulr_cg = new(); clmulr_cg.set_inst_name("obj_clmulr");
