///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
// 
// Copyright (C) 2024 Harvey Mudd College, 10x Engineers, UET Lahore, Habib University
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
////////////////////////////////////////////////////////////////////////////////////////////////

    cbo_inval_cg = new(); cbo_inval_cg.set_inst_name("obj_cbo_inval");
    cbo_clean_cg = new(); cbo_clean_cg.set_inst_name("obj_cbo_clean");
    cbo_flush_cg = new(); cbo_flush_cg.set_inst_name("obj_cbo_flush");